.include TSMC_180nm.txt


.param SUPPLY = 1.8

.global gnd

Vdd vdd gnd 'SUPPLY'

V_in_a node_in gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)

* SPICE3 file created from not.ext - technology: scmos

.option scale=0.09u

M1000 node_out node_in gnd Gnd CMOSN w=14 l=4
+  ad=336 pd=76 as=336 ps=76
M1001 node_out node_in vdd vdd CMOSP w=10 l=4
+  ad=240 pd=68 as=240 ps=68
C0 gnd node_in 0.05fF
C1 vdd node_out 0.03fF
C2 vdd vdd 0.02fF
C3 node_in vdd 0.05fF
C4 vdd node_in 0.11fF
C5 gnd Gnd 0.30fF
C6 node_out Gnd 0.08fF
C7 vdd Gnd 0.25fF
C8 node_in Gnd 0.43fF
C9 vdd Gnd 1.66fF

C10 node_out gnd 75fF
.tran 1n 800n

.measure tran trise 
+ TRIG v(node_in) VAL = 'SUPPLY/2' RISE =1
+ TARG v(node_out) VAL = 'SUPPLY/2' FALL =1 

.measure tran tfall 
+ TRIG v(node_in) VAL = 'SUPPLY/2' FALL =1 
+ TARG v(node_out) VAL = 'SUPPLY/2' RISE=1

.measure tran tpd param = '(trise + tfall)/2' goal = 0

.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(node_in) v(node_out)+2
hardcopy image.ps v(node_in)  v(node_out)+2
.end
.endc