magic
tech scmos
timestamp 1700146955
<< nwell >>
rect -280 176 -92 215
rect -53 176 47 206
rect 120 162 190 178
rect -37 37 63 67
rect -270 -80 -82 -41
<< ntransistor >>
rect -38 130 -34 139
rect -6 130 -2 139
rect 28 130 32 139
rect 135 127 137 131
rect 153 127 155 131
rect 172 127 174 131
rect -265 118 -262 125
rect -236 118 -234 125
rect -205 118 -202 125
rect -176 118 -173 125
rect -147 118 -144 125
rect -117 118 -114 125
rect -22 -9 -18 0
rect 10 -9 14 0
rect 44 -9 48 0
rect -255 -138 -252 -131
rect -226 -138 -224 -131
rect -195 -138 -192 -131
rect -166 -138 -163 -131
rect -137 -138 -134 -131
rect -107 -138 -104 -131
<< ptransistor >>
rect -265 190 -262 197
rect -236 190 -234 197
rect -205 190 -202 197
rect -176 190 -173 197
rect -147 190 -144 197
rect -117 190 -114 197
rect -38 188 -34 197
rect -6 188 -2 197
rect 28 188 32 197
rect 135 168 137 172
rect 153 168 155 172
rect 172 168 174 172
rect -22 49 -18 58
rect 10 49 14 58
rect 44 49 48 58
rect -255 -66 -252 -59
rect -226 -66 -224 -59
rect -195 -66 -192 -59
rect -166 -66 -163 -59
rect -137 -66 -134 -59
rect -107 -66 -104 -59
<< ndiffusion >>
rect -42 134 -38 139
rect -47 130 -38 134
rect -34 134 -28 139
rect -34 130 -23 134
rect -11 134 -6 139
rect -16 130 -6 134
rect -2 134 3 139
rect -2 130 8 134
rect 22 134 28 139
rect 17 130 28 134
rect 32 134 36 139
rect 32 130 41 134
rect 133 127 135 131
rect 137 127 139 131
rect 151 127 153 131
rect 155 127 157 131
rect 170 127 172 131
rect 174 127 176 131
rect -270 121 -265 125
rect -274 118 -265 121
rect -262 121 -253 125
rect -262 118 -249 121
rect -241 121 -236 125
rect -245 118 -236 121
rect -234 121 -224 125
rect -234 118 -220 121
rect -212 121 -205 125
rect -216 118 -205 121
rect -202 121 -195 125
rect -202 118 -191 121
rect -183 121 -176 125
rect -187 118 -176 121
rect -173 121 -166 125
rect -173 118 -162 121
rect -154 121 -147 125
rect -158 118 -147 121
rect -144 121 -137 125
rect -144 118 -133 121
rect -125 121 -117 125
rect -129 118 -117 121
rect -114 121 -108 125
rect -114 118 -104 121
rect -26 -5 -22 0
rect -31 -9 -22 -5
rect -18 -5 -12 0
rect -18 -9 -7 -5
rect 5 -5 10 0
rect 0 -9 10 -5
rect 14 -5 19 0
rect 14 -9 24 -5
rect 38 -5 44 0
rect 33 -9 44 -5
rect 48 -5 52 0
rect 48 -9 57 -5
rect -260 -135 -255 -131
rect -264 -138 -255 -135
rect -252 -135 -243 -131
rect -252 -138 -239 -135
rect -231 -135 -226 -131
rect -235 -138 -226 -135
rect -224 -135 -214 -131
rect -224 -138 -210 -135
rect -202 -135 -195 -131
rect -206 -138 -195 -135
rect -192 -135 -185 -131
rect -192 -138 -181 -135
rect -173 -135 -166 -131
rect -177 -138 -166 -135
rect -163 -135 -156 -131
rect -163 -138 -152 -135
rect -144 -135 -137 -131
rect -148 -138 -137 -135
rect -134 -135 -127 -131
rect -134 -138 -123 -135
rect -115 -135 -107 -131
rect -119 -138 -107 -135
rect -104 -135 -98 -131
rect -104 -138 -94 -135
<< pdiffusion >>
rect -270 193 -265 197
rect -274 190 -265 193
rect -262 193 -253 197
rect -262 190 -249 193
rect -241 193 -236 197
rect -245 190 -236 193
rect -234 193 -224 197
rect -234 190 -220 193
rect -212 193 -205 197
rect -216 190 -205 193
rect -202 193 -195 197
rect -202 190 -191 193
rect -183 193 -176 197
rect -187 190 -176 193
rect -173 193 -166 197
rect -173 190 -162 193
rect -154 193 -147 197
rect -158 190 -147 193
rect -144 193 -137 197
rect -144 190 -133 193
rect -125 193 -117 197
rect -129 190 -117 193
rect -114 193 -108 197
rect -114 190 -104 193
rect -42 192 -38 197
rect -47 188 -38 192
rect -34 192 -28 197
rect -34 188 -23 192
rect -11 192 -6 197
rect -16 188 -6 192
rect -2 192 3 197
rect -2 188 8 192
rect 22 192 28 197
rect 17 188 28 192
rect 32 192 36 197
rect 32 188 41 192
rect 133 168 135 172
rect 137 168 139 172
rect 151 168 153 172
rect 155 168 157 172
rect 170 168 172 172
rect 174 168 176 172
rect -26 53 -22 58
rect -31 49 -22 53
rect -18 53 -12 58
rect -18 49 -7 53
rect 5 53 10 58
rect 0 49 10 53
rect 14 53 19 58
rect 14 49 24 53
rect 38 53 44 58
rect 33 49 44 53
rect 48 53 52 58
rect 48 49 57 53
rect -260 -63 -255 -59
rect -264 -66 -255 -63
rect -252 -63 -243 -59
rect -252 -66 -239 -63
rect -231 -63 -226 -59
rect -235 -66 -226 -63
rect -224 -63 -214 -59
rect -224 -66 -210 -63
rect -202 -63 -195 -59
rect -206 -66 -195 -63
rect -192 -63 -185 -59
rect -192 -66 -181 -63
rect -173 -63 -166 -59
rect -177 -66 -166 -63
rect -163 -63 -156 -59
rect -163 -66 -152 -63
rect -144 -63 -137 -59
rect -148 -66 -137 -63
rect -134 -63 -127 -59
rect -134 -66 -123 -63
rect -115 -63 -107 -59
rect -119 -66 -107 -63
rect -104 -63 -98 -59
rect -104 -66 -94 -63
<< ndcontact >>
rect -47 134 -42 139
rect -28 134 -23 139
rect -16 134 -11 139
rect 3 134 8 139
rect 17 134 22 139
rect 36 134 41 139
rect 129 127 133 131
rect 139 127 143 131
rect 147 127 151 131
rect 157 127 161 131
rect 166 127 170 131
rect 176 127 180 131
rect -274 121 -270 125
rect -253 121 -249 125
rect -245 121 -241 125
rect -224 121 -220 125
rect -216 121 -212 125
rect -195 121 -191 125
rect -187 121 -183 125
rect -166 121 -162 125
rect -158 121 -154 125
rect -137 121 -133 125
rect -129 121 -125 125
rect -108 121 -104 125
rect -31 -5 -26 0
rect -12 -5 -7 0
rect 0 -5 5 0
rect 19 -5 24 0
rect 33 -5 38 0
rect 52 -5 57 0
rect -264 -135 -260 -131
rect -243 -135 -239 -131
rect -235 -135 -231 -131
rect -214 -135 -210 -131
rect -206 -135 -202 -131
rect -185 -135 -181 -131
rect -177 -135 -173 -131
rect -156 -135 -152 -131
rect -148 -135 -144 -131
rect -127 -135 -123 -131
rect -119 -135 -115 -131
rect -98 -135 -94 -131
<< pdcontact >>
rect -274 193 -270 197
rect -253 193 -249 197
rect -245 193 -241 197
rect -224 193 -220 197
rect -216 193 -212 197
rect -195 193 -191 197
rect -187 193 -183 197
rect -166 193 -162 197
rect -158 193 -154 197
rect -137 193 -133 197
rect -129 193 -125 197
rect -108 193 -104 197
rect -47 192 -42 197
rect -28 192 -23 197
rect -16 192 -11 197
rect 3 192 8 197
rect 17 192 22 197
rect 36 192 41 197
rect 129 168 133 172
rect 139 168 143 172
rect 147 168 151 172
rect 157 168 161 172
rect 166 168 170 172
rect 176 168 180 172
rect -31 53 -26 58
rect -12 53 -7 58
rect 0 53 5 58
rect 19 53 24 58
rect 33 53 38 58
rect 52 53 57 58
rect -264 -63 -260 -59
rect -243 -63 -239 -59
rect -235 -63 -231 -59
rect -214 -63 -210 -59
rect -206 -63 -202 -59
rect -185 -63 -181 -59
rect -177 -63 -173 -59
rect -156 -63 -152 -59
rect -148 -63 -144 -59
rect -127 -63 -123 -59
rect -119 -63 -115 -59
rect -98 -63 -94 -59
<< polysilicon >>
rect -265 203 -202 205
rect -265 197 -262 203
rect -236 197 -234 200
rect -205 197 -202 203
rect -176 197 -173 201
rect -147 197 -144 201
rect -117 197 -114 201
rect -38 197 -34 203
rect -6 197 -2 201
rect 28 197 32 201
rect -265 125 -262 190
rect -236 125 -234 190
rect -205 125 -202 190
rect -176 125 -173 190
rect -154 163 -151 168
rect -147 125 -144 190
rect -117 125 -114 190
rect -38 154 -34 188
rect -37 149 -34 154
rect -38 139 -34 149
rect -6 139 -2 188
rect 28 139 32 188
rect 135 172 137 175
rect 153 172 155 175
rect 172 172 174 175
rect 135 145 137 168
rect 153 147 155 168
rect 172 148 174 168
rect 136 141 137 145
rect 154 143 155 147
rect 173 144 174 148
rect 135 131 137 141
rect 153 131 155 143
rect 172 131 174 144
rect -38 127 -34 130
rect -6 127 -2 130
rect 28 127 32 130
rect 135 124 137 127
rect 153 124 155 127
rect 172 124 174 127
rect -265 113 -262 118
rect -236 106 -234 118
rect -205 115 -202 118
rect -176 106 -173 118
rect -147 113 -144 118
rect -117 113 -114 118
rect -236 103 -173 106
rect -22 58 -18 64
rect 10 58 14 62
rect 44 58 48 62
rect -22 15 -18 49
rect -21 10 -18 15
rect -22 0 -18 10
rect 10 0 14 49
rect 44 0 48 49
rect -22 -12 -18 -9
rect 10 -12 14 -9
rect 44 -12 48 -9
rect -255 -53 -192 -51
rect -255 -59 -252 -53
rect -226 -59 -224 -56
rect -195 -59 -192 -53
rect -166 -59 -163 -55
rect -137 -59 -134 -55
rect -107 -59 -104 -55
rect -255 -131 -252 -66
rect -226 -131 -224 -66
rect -195 -131 -192 -66
rect -166 -131 -163 -66
rect -144 -93 -141 -88
rect -137 -131 -134 -66
rect -107 -131 -104 -66
rect -255 -143 -252 -138
rect -226 -150 -224 -138
rect -195 -141 -192 -138
rect -166 -150 -163 -138
rect -137 -143 -134 -138
rect -107 -143 -104 -138
rect -226 -153 -163 -150
<< polycontact >>
rect -270 154 -265 159
rect -241 153 -236 158
rect -151 163 -147 168
rect -122 136 -117 142
rect -41 149 -37 154
rect -10 149 -6 154
rect 22 162 28 168
rect 132 141 136 145
rect 150 143 154 147
rect 169 144 173 148
rect -25 10 -21 15
rect 6 10 10 15
rect 38 23 44 29
rect -260 -102 -255 -97
rect -231 -103 -226 -98
rect -141 -93 -137 -88
rect -112 -120 -107 -114
<< metal1 >>
rect -337 216 -67 222
rect -337 215 -264 216
rect -337 -26 -323 215
rect -274 197 -270 215
rect -245 197 -241 216
rect -216 197 -212 216
rect -187 197 -183 216
rect -72 213 -67 216
rect -72 206 201 213
rect -166 202 -125 206
rect -166 197 -162 202
rect -158 197 -154 202
rect -129 197 -125 202
rect -47 197 -42 206
rect -16 197 -11 206
rect 17 197 22 206
rect -253 169 -249 193
rect -253 165 -233 169
rect -272 154 -270 159
rect -253 125 -249 165
rect -224 142 -220 193
rect -195 186 -191 193
rect -166 186 -162 193
rect -195 183 -162 186
rect -137 186 -133 193
rect -108 186 -104 193
rect -137 183 -104 186
rect -159 164 -151 168
rect -154 163 -151 164
rect -108 160 -104 183
rect -28 168 -23 192
rect 3 168 8 192
rect -28 162 22 168
rect -108 157 -100 160
rect -108 152 -66 157
rect -108 150 -100 152
rect -224 137 -122 142
rect -224 125 -220 137
rect -126 136 -122 137
rect -108 133 -104 150
rect -166 125 -162 126
rect -108 125 -104 128
rect -191 121 -187 125
rect -133 121 -129 125
rect -274 117 -270 121
rect -245 117 -241 121
rect -216 117 -212 121
rect -158 117 -154 121
rect -302 110 -96 117
rect -302 -139 -290 110
rect -73 15 -66 152
rect -42 149 -41 154
rect -11 149 -10 154
rect 3 139 8 162
rect 36 139 41 192
rect 195 183 201 206
rect 115 178 201 183
rect 129 172 133 178
rect 166 172 170 178
rect 143 168 147 172
rect 157 148 161 168
rect 176 151 180 168
rect -23 134 -16 139
rect 110 141 132 145
rect 149 143 150 147
rect 157 144 169 148
rect 176 147 185 151
rect 110 140 131 141
rect -47 130 -42 134
rect 17 130 22 134
rect -53 129 48 130
rect -46 123 48 129
rect -38 67 91 74
rect -31 58 -26 67
rect 0 58 5 67
rect 33 58 38 67
rect -12 29 -7 53
rect 19 29 24 53
rect -12 23 38 29
rect 52 26 57 53
rect 110 26 117 140
rect 157 139 161 144
rect 139 136 161 139
rect 139 131 143 136
rect 157 131 161 136
rect 176 131 180 147
rect 129 124 133 127
rect 147 124 151 127
rect 166 124 170 127
rect 125 123 189 124
rect 134 121 189 123
rect 194 74 201 178
rect 157 67 201 74
rect -73 10 -25 15
rect 3 10 6 15
rect -262 -39 -82 -33
rect -270 -40 -82 -39
rect -264 -59 -260 -40
rect -235 -59 -231 -40
rect -206 -59 -202 -40
rect -177 -59 -173 -40
rect -156 -54 -115 -50
rect -156 -59 -152 -54
rect -148 -59 -144 -54
rect -119 -59 -115 -54
rect -263 -102 -260 -97
rect -243 -131 -239 -63
rect -214 -114 -210 -63
rect -185 -70 -181 -63
rect -156 -70 -152 -63
rect -185 -73 -152 -70
rect -127 -70 -123 -63
rect -98 -70 -94 -63
rect -127 -73 -94 -70
rect -149 -92 -141 -88
rect -144 -93 -141 -92
rect -98 -96 -94 -73
rect -98 -106 -90 -96
rect -214 -119 -112 -114
rect -214 -131 -210 -119
rect -116 -120 -112 -119
rect -98 -123 -94 -106
rect -156 -131 -152 -130
rect -98 -131 -94 -128
rect -181 -135 -177 -131
rect -123 -135 -119 -131
rect -264 -139 -260 -135
rect -235 -139 -231 -135
rect -206 -139 -202 -135
rect -148 -139 -144 -135
rect -302 -146 -79 -139
rect -302 -204 -290 -146
rect -73 -167 -66 10
rect 19 0 24 23
rect 52 21 117 26
rect 52 0 57 21
rect -7 -5 0 0
rect -31 -9 -26 -5
rect 33 -9 38 -5
rect -229 -174 -66 -167
rect -37 -16 70 -9
rect -37 -204 -23 -16
rect -302 -213 -23 -204
<< m2contact >>
rect -277 154 -272 159
rect -233 164 -227 169
rect -246 153 -241 158
rect -164 164 -159 169
rect -166 126 -161 131
rect -109 128 -104 133
rect -337 -40 -323 -26
rect -96 110 -87 118
rect -47 149 -42 154
rect -16 149 -11 154
rect 41 160 49 165
rect 144 143 149 148
rect -55 121 -46 129
rect 48 122 57 130
rect 91 67 101 74
rect 125 115 134 123
rect 148 67 157 74
rect -3 10 3 16
rect -270 -39 -262 -32
rect -269 -102 -263 -96
rect -239 -92 -233 -87
rect -236 -103 -231 -98
rect -154 -92 -149 -87
rect -156 -130 -151 -125
rect -99 -128 -94 -123
rect -234 -174 -229 -167
<< metal2 >>
rect -246 225 -12 228
rect -277 149 -272 154
rect -246 158 -242 225
rect -227 164 -164 168
rect -16 154 -12 225
rect 78 189 149 193
rect 78 165 82 189
rect 49 160 82 165
rect -128 149 -47 153
rect -277 146 -124 149
rect 144 148 149 189
rect -161 128 -109 131
rect -55 116 -46 121
rect -87 110 -46 116
rect -96 109 -46 110
rect 49 111 56 122
rect 125 111 134 115
rect 49 106 134 111
rect 101 67 148 74
rect -323 -39 -270 -34
rect -323 -40 -264 -39
rect -233 -92 -154 -88
rect -269 -186 -263 -102
rect -234 -167 -231 -103
rect -151 -128 -99 -125
rect -3 -186 3 10
rect -269 -190 3 -186
<< labels >>
rlabel metal1 -272 156 -272 156 1 node_a
rlabel m2contact -243 154 -243 154 1 node_b
rlabel metal1 -215 115 -215 115 1 gnd
rlabel metal1 -105 155 -105 155 1 node_y1
rlabel metal1 39 162 39 162 1 node_y2
rlabel metal1 181 148 181 148 1 node_c
rlabel m2contact -264 -101 -264 -101 1 node_cin
rlabel metal1 -94 -100 -94 -100 1 node_s
rlabel metal1 -234 219 -234 219 5 vdd
rlabel metal1 54 22 54 22 1 node_y3
<< end >>
