magic
tech scmos
timestamp 1700174420
<< nwell >>
rect -341 1125 -266 1147
rect -71 1120 4 1142
rect 184 1126 259 1148
rect 452 1126 527 1148
rect 1011 971 1189 1006
rect -195 914 80 955
rect 187 914 462 955
rect 569 914 844 955
rect -373 852 -273 882
rect -357 597 -153 629
rect -358 350 -154 382
rect -4 294 271 335
rect -354 124 -150 156
rect -357 -83 -153 -51
<< ntransistor >>
rect -307 1089 -303 1103
rect -37 1084 -33 1098
rect 218 1090 222 1104
rect 486 1090 490 1104
rect 1030 903 1034 912
rect 1065 903 1069 912
rect 1098 903 1102 912
rect 1131 903 1135 912
rect 1164 903 1168 912
rect -173 830 -169 841
rect -127 830 -123 841
rect -82 830 -78 841
rect -39 830 -35 841
rect 6 830 10 841
rect 49 830 53 841
rect 209 830 213 841
rect 255 830 259 841
rect 300 830 304 841
rect 343 830 347 841
rect 388 830 392 841
rect 431 830 435 841
rect 591 830 595 841
rect 637 830 641 841
rect 682 830 686 841
rect 725 830 729 841
rect 770 830 774 841
rect 813 830 817 841
rect -358 806 -354 815
rect -326 806 -322 815
rect -292 806 -288 815
rect -341 522 -338 528
rect -306 522 -303 528
rect -271 522 -268 528
rect -239 522 -236 528
rect -208 522 -205 528
rect -175 522 -172 528
rect -342 275 -339 281
rect -307 275 -304 281
rect -272 275 -269 281
rect -240 275 -237 281
rect -209 275 -206 281
rect -176 275 -173 281
rect 18 210 22 221
rect 64 210 68 221
rect 109 210 113 221
rect 152 210 156 221
rect 197 210 201 221
rect 240 210 244 221
rect -338 49 -335 55
rect -303 49 -300 55
rect -268 49 -265 55
rect -236 49 -233 55
rect -205 49 -202 55
rect -172 49 -169 55
rect -341 -158 -338 -152
rect -306 -158 -303 -152
rect -271 -158 -268 -152
rect -239 -158 -236 -152
rect -208 -158 -205 -152
rect -175 -158 -172 -152
<< ptransistor >>
rect -307 1131 -303 1141
rect -37 1126 -33 1136
rect 218 1132 222 1142
rect 486 1132 490 1142
rect 1030 985 1034 994
rect 1065 985 1069 994
rect 1098 985 1102 994
rect 1131 985 1135 994
rect 1164 985 1168 994
rect -173 933 -169 944
rect -127 933 -123 944
rect -82 933 -78 944
rect -39 933 -35 944
rect 6 933 10 944
rect 49 933 53 944
rect 209 933 213 944
rect 255 933 259 944
rect 300 933 304 944
rect 343 933 347 944
rect 388 933 392 944
rect 431 933 435 944
rect 591 933 595 944
rect 637 933 641 944
rect 682 933 686 944
rect 725 933 729 944
rect 770 933 774 944
rect 813 933 817 944
rect -358 864 -354 873
rect -326 864 -322 873
rect -292 864 -288 873
rect -341 611 -338 617
rect -306 611 -303 617
rect -271 611 -268 617
rect -239 611 -236 617
rect -208 611 -205 617
rect -175 611 -172 617
rect -342 364 -339 370
rect -307 364 -304 370
rect -272 364 -269 370
rect -240 364 -237 370
rect -209 364 -206 370
rect -176 364 -173 370
rect 18 313 22 324
rect 64 313 68 324
rect 109 313 113 324
rect 152 313 156 324
rect 197 313 201 324
rect 240 313 244 324
rect -338 138 -335 144
rect -303 138 -300 144
rect -268 138 -265 144
rect -236 138 -233 144
rect -205 138 -202 144
rect -172 138 -169 144
rect -341 -69 -338 -63
rect -306 -69 -303 -63
rect -271 -69 -268 -63
rect -239 -69 -236 -63
rect -208 -69 -205 -63
rect -175 -69 -172 -63
<< ndiffusion >>
rect -327 1099 -307 1103
rect -331 1089 -307 1099
rect -303 1099 -283 1103
rect -303 1089 -279 1099
rect 198 1100 218 1104
rect -57 1094 -37 1098
rect -61 1084 -37 1094
rect -33 1094 -13 1098
rect -33 1084 -9 1094
rect 194 1090 218 1100
rect 222 1100 242 1104
rect 222 1090 246 1100
rect 466 1100 486 1104
rect 462 1090 486 1100
rect 490 1100 510 1104
rect 490 1090 514 1100
rect 1022 908 1030 912
rect 1018 903 1030 908
rect 1034 908 1043 912
rect 1034 903 1047 908
rect 1056 908 1065 912
rect 1052 903 1065 908
rect 1069 908 1077 912
rect 1069 903 1081 908
rect 1089 908 1098 912
rect 1085 903 1098 908
rect 1102 908 1110 912
rect 1102 903 1114 908
rect 1122 908 1131 912
rect 1118 903 1131 908
rect 1135 908 1143 912
rect 1135 903 1147 908
rect 1155 908 1164 912
rect 1151 903 1164 908
rect 1168 908 1176 912
rect 1168 903 1180 908
rect -185 837 -173 841
rect -189 830 -173 837
rect -169 837 -153 841
rect -169 830 -149 837
rect -141 837 -127 841
rect -145 830 -127 837
rect -123 837 -109 841
rect -123 830 -105 837
rect -97 837 -82 841
rect -101 830 -82 837
rect -78 837 -65 841
rect -78 830 -61 837
rect -53 837 -39 841
rect -57 830 -39 837
rect -35 837 -21 841
rect -35 830 -17 837
rect -9 837 6 841
rect -13 830 6 837
rect 10 837 23 841
rect 10 830 27 837
rect 35 837 49 841
rect 31 830 49 837
rect 53 837 67 841
rect 53 830 71 837
rect 197 837 209 841
rect 193 830 209 837
rect 213 837 229 841
rect 213 830 233 837
rect 241 837 255 841
rect 237 830 255 837
rect 259 837 273 841
rect 259 830 277 837
rect 285 837 300 841
rect 281 830 300 837
rect 304 837 317 841
rect 304 830 321 837
rect 329 837 343 841
rect 325 830 343 837
rect 347 837 361 841
rect 347 830 365 837
rect 373 837 388 841
rect 369 830 388 837
rect 392 837 405 841
rect 392 830 409 837
rect 417 837 431 841
rect 413 830 431 837
rect 435 837 449 841
rect 435 830 453 837
rect 579 837 591 841
rect 575 830 591 837
rect 595 837 611 841
rect 595 830 615 837
rect 623 837 637 841
rect 619 830 637 837
rect 641 837 655 841
rect 641 830 659 837
rect 667 837 682 841
rect 663 830 682 837
rect 686 837 699 841
rect 686 830 703 837
rect 711 837 725 841
rect 707 830 725 837
rect 729 837 743 841
rect 729 830 747 837
rect 755 837 770 841
rect 751 830 770 837
rect 774 837 787 841
rect 774 830 791 837
rect 799 837 813 841
rect 795 830 813 837
rect 817 837 831 841
rect 817 830 835 837
rect -362 810 -358 815
rect -367 806 -358 810
rect -354 810 -348 815
rect -354 806 -343 810
rect -331 810 -326 815
rect -336 806 -326 810
rect -322 810 -317 815
rect -322 806 -312 810
rect -298 810 -292 815
rect -303 806 -292 810
rect -288 810 -284 815
rect -288 806 -279 810
rect -347 524 -341 528
rect -351 522 -341 524
rect -338 524 -328 528
rect -338 522 -324 524
rect -313 524 -306 528
rect -317 522 -306 524
rect -303 524 -294 528
rect -303 522 -290 524
rect -280 524 -271 528
rect -284 522 -271 524
rect -268 524 -261 528
rect -268 522 -257 524
rect -248 524 -239 528
rect -252 522 -239 524
rect -236 524 -229 528
rect -236 522 -225 524
rect -216 524 -208 528
rect -220 522 -208 524
rect -205 524 -197 528
rect -205 522 -193 524
rect -184 524 -175 528
rect -188 522 -175 524
rect -172 524 -165 528
rect -172 522 -161 524
rect -348 277 -342 281
rect -352 275 -342 277
rect -339 277 -329 281
rect -339 275 -325 277
rect -314 277 -307 281
rect -318 275 -307 277
rect -304 277 -295 281
rect -304 275 -291 277
rect -281 277 -272 281
rect -285 275 -272 277
rect -269 277 -262 281
rect -269 275 -258 277
rect -249 277 -240 281
rect -253 275 -240 277
rect -237 277 -230 281
rect -237 275 -226 277
rect -217 277 -209 281
rect -221 275 -209 277
rect -206 277 -198 281
rect -206 275 -194 277
rect -185 277 -176 281
rect -189 275 -176 277
rect -173 277 -166 281
rect -173 275 -162 277
rect 6 217 18 221
rect 2 210 18 217
rect 22 217 38 221
rect 22 210 42 217
rect 50 217 64 221
rect 46 210 64 217
rect 68 217 82 221
rect 68 210 86 217
rect 94 217 109 221
rect 90 210 109 217
rect 113 217 126 221
rect 113 210 130 217
rect 138 217 152 221
rect 134 210 152 217
rect 156 217 170 221
rect 156 210 174 217
rect 182 217 197 221
rect 178 210 197 217
rect 201 217 214 221
rect 201 210 218 217
rect 226 217 240 221
rect 222 210 240 217
rect 244 217 258 221
rect 244 210 262 217
rect -344 51 -338 55
rect -348 49 -338 51
rect -335 51 -325 55
rect -335 49 -321 51
rect -310 51 -303 55
rect -314 49 -303 51
rect -300 51 -291 55
rect -300 49 -287 51
rect -277 51 -268 55
rect -281 49 -268 51
rect -265 51 -258 55
rect -265 49 -254 51
rect -245 51 -236 55
rect -249 49 -236 51
rect -233 51 -226 55
rect -233 49 -222 51
rect -213 51 -205 55
rect -217 49 -205 51
rect -202 51 -194 55
rect -202 49 -190 51
rect -181 51 -172 55
rect -185 49 -172 51
rect -169 51 -162 55
rect -169 49 -158 51
rect -347 -156 -341 -152
rect -351 -158 -341 -156
rect -338 -156 -328 -152
rect -338 -158 -324 -156
rect -313 -156 -306 -152
rect -317 -158 -306 -156
rect -303 -156 -294 -152
rect -303 -158 -290 -156
rect -280 -156 -271 -152
rect -284 -158 -271 -156
rect -268 -156 -261 -152
rect -268 -158 -257 -156
rect -248 -156 -239 -152
rect -252 -158 -239 -156
rect -236 -156 -229 -152
rect -236 -158 -225 -156
rect -216 -156 -208 -152
rect -220 -158 -208 -156
rect -205 -156 -197 -152
rect -205 -158 -193 -156
rect -184 -156 -175 -152
rect -188 -158 -175 -156
rect -172 -156 -165 -152
rect -172 -158 -161 -156
<< pdiffusion >>
rect -327 1137 -307 1141
rect -331 1131 -307 1137
rect -303 1137 -283 1141
rect -303 1131 -279 1137
rect 198 1138 218 1142
rect -57 1132 -37 1136
rect -61 1126 -37 1132
rect -33 1132 -13 1136
rect 194 1132 218 1138
rect 222 1138 242 1142
rect 222 1132 246 1138
rect 466 1138 486 1142
rect 462 1132 486 1138
rect 490 1138 510 1142
rect 490 1132 514 1138
rect -33 1126 -9 1132
rect 1022 990 1030 994
rect 1018 985 1030 990
rect 1034 990 1043 994
rect 1034 985 1047 990
rect 1056 990 1065 994
rect 1052 985 1065 990
rect 1069 990 1077 994
rect 1069 985 1081 990
rect 1089 990 1098 994
rect 1085 985 1098 990
rect 1102 990 1110 994
rect 1102 985 1114 990
rect 1122 990 1131 994
rect 1118 985 1131 990
rect 1135 990 1143 994
rect 1135 985 1147 990
rect 1155 990 1164 994
rect 1151 985 1164 990
rect 1168 990 1176 994
rect 1168 985 1180 990
rect -185 940 -173 944
rect -189 933 -173 940
rect -169 940 -153 944
rect -169 933 -149 940
rect -141 940 -127 944
rect -145 933 -127 940
rect -123 940 -109 944
rect -123 933 -105 940
rect -97 940 -82 944
rect -101 933 -82 940
rect -78 940 -65 944
rect -78 933 -61 940
rect -53 940 -39 944
rect -57 933 -39 940
rect -35 940 -21 944
rect -35 933 -17 940
rect -9 940 6 944
rect -13 933 6 940
rect 10 940 23 944
rect 10 933 27 940
rect 35 940 49 944
rect 31 933 49 940
rect 53 940 67 944
rect 53 933 71 940
rect 197 940 209 944
rect 193 933 209 940
rect 213 940 229 944
rect 213 933 233 940
rect 241 940 255 944
rect 237 933 255 940
rect 259 940 273 944
rect 259 933 277 940
rect 285 940 300 944
rect 281 933 300 940
rect 304 940 317 944
rect 304 933 321 940
rect 329 940 343 944
rect 325 933 343 940
rect 347 940 361 944
rect 347 933 365 940
rect 373 940 388 944
rect 369 933 388 940
rect 392 940 405 944
rect 392 933 409 940
rect 417 940 431 944
rect 413 933 431 940
rect 435 940 449 944
rect 435 933 453 940
rect 579 940 591 944
rect 575 933 591 940
rect 595 940 611 944
rect 595 933 615 940
rect 623 940 637 944
rect 619 933 637 940
rect 641 940 655 944
rect 641 933 659 940
rect 667 940 682 944
rect 663 933 682 940
rect 686 940 699 944
rect 686 933 703 940
rect 711 940 725 944
rect 707 933 725 940
rect 729 940 743 944
rect 729 933 747 940
rect 755 940 770 944
rect 751 933 770 940
rect 774 940 787 944
rect 774 933 791 940
rect 799 940 813 944
rect 795 933 813 940
rect 817 940 831 944
rect 817 933 835 940
rect -362 868 -358 873
rect -367 864 -358 868
rect -354 868 -348 873
rect -354 864 -343 868
rect -331 868 -326 873
rect -336 864 -326 868
rect -322 868 -317 873
rect -322 864 -312 868
rect -298 868 -292 873
rect -303 864 -292 868
rect -288 868 -284 873
rect -288 864 -279 868
rect -347 613 -341 617
rect -351 611 -341 613
rect -338 613 -328 617
rect -338 611 -324 613
rect -313 613 -306 617
rect -317 611 -306 613
rect -303 613 -294 617
rect -303 611 -290 613
rect -280 613 -271 617
rect -284 611 -271 613
rect -268 613 -261 617
rect -268 611 -257 613
rect -248 613 -239 617
rect -252 611 -239 613
rect -236 613 -229 617
rect -236 611 -225 613
rect -216 613 -208 617
rect -220 611 -208 613
rect -205 613 -197 617
rect -205 611 -193 613
rect -184 613 -175 617
rect -188 611 -175 613
rect -172 613 -165 617
rect -172 611 -161 613
rect -348 366 -342 370
rect -352 364 -342 366
rect -339 366 -329 370
rect -339 364 -325 366
rect -314 366 -307 370
rect -318 364 -307 366
rect -304 366 -295 370
rect -304 364 -291 366
rect -281 366 -272 370
rect -285 364 -272 366
rect -269 366 -262 370
rect -269 364 -258 366
rect -249 366 -240 370
rect -253 364 -240 366
rect -237 366 -230 370
rect -237 364 -226 366
rect -217 366 -209 370
rect -221 364 -209 366
rect -206 366 -198 370
rect -206 364 -194 366
rect -185 366 -176 370
rect -189 364 -176 366
rect -173 366 -166 370
rect -173 364 -162 366
rect 6 320 18 324
rect 2 313 18 320
rect 22 320 38 324
rect 22 313 42 320
rect 50 320 64 324
rect 46 313 64 320
rect 68 320 82 324
rect 68 313 86 320
rect 94 320 109 324
rect 90 313 109 320
rect 113 320 126 324
rect 113 313 130 320
rect 138 320 152 324
rect 134 313 152 320
rect 156 320 170 324
rect 156 313 174 320
rect 182 320 197 324
rect 178 313 197 320
rect 201 320 214 324
rect 201 313 218 320
rect 226 320 240 324
rect 222 313 240 320
rect 244 320 258 324
rect 244 313 262 320
rect -344 140 -338 144
rect -348 138 -338 140
rect -335 140 -325 144
rect -335 138 -321 140
rect -310 140 -303 144
rect -314 138 -303 140
rect -300 140 -291 144
rect -300 138 -287 140
rect -277 140 -268 144
rect -281 138 -268 140
rect -265 140 -258 144
rect -265 138 -254 140
rect -245 140 -236 144
rect -249 138 -236 140
rect -233 140 -226 144
rect -233 138 -222 140
rect -213 140 -205 144
rect -217 138 -205 140
rect -202 140 -194 144
rect -202 138 -190 140
rect -181 140 -172 144
rect -185 138 -172 140
rect -169 140 -162 144
rect -169 138 -158 140
rect -347 -67 -341 -63
rect -351 -69 -341 -67
rect -338 -67 -328 -63
rect -338 -69 -324 -67
rect -313 -67 -306 -63
rect -317 -69 -306 -67
rect -303 -67 -294 -63
rect -303 -69 -290 -67
rect -280 -67 -271 -63
rect -284 -69 -271 -67
rect -268 -67 -261 -63
rect -268 -69 -257 -67
rect -248 -67 -239 -63
rect -252 -69 -239 -67
rect -236 -67 -229 -63
rect -236 -69 -225 -67
rect -216 -67 -208 -63
rect -220 -69 -208 -67
rect -205 -67 -197 -63
rect -205 -69 -193 -67
rect -184 -67 -175 -63
rect -188 -69 -175 -67
rect -172 -67 -165 -63
rect -172 -69 -161 -67
<< ndcontact >>
rect -331 1099 -327 1103
rect -283 1099 -279 1103
rect 194 1100 198 1104
rect -61 1094 -57 1098
rect -13 1094 -9 1098
rect 242 1100 246 1104
rect 462 1100 466 1104
rect 510 1100 514 1104
rect 1018 908 1022 912
rect 1043 908 1047 912
rect 1052 908 1056 912
rect 1077 908 1081 912
rect 1085 908 1089 912
rect 1110 908 1114 912
rect 1118 908 1122 912
rect 1143 908 1147 912
rect 1151 908 1155 912
rect 1176 908 1180 912
rect -189 837 -185 841
rect -153 837 -149 841
rect -145 837 -141 841
rect -109 837 -105 841
rect -101 837 -97 841
rect -65 837 -61 841
rect -57 837 -53 841
rect -21 837 -17 841
rect -13 837 -9 841
rect 23 837 27 841
rect 31 837 35 841
rect 67 837 71 841
rect 193 837 197 841
rect 229 837 233 841
rect 237 837 241 841
rect 273 837 277 841
rect 281 837 285 841
rect 317 837 321 841
rect 325 837 329 841
rect 361 837 365 841
rect 369 837 373 841
rect 405 837 409 841
rect 413 837 417 841
rect 449 837 453 841
rect 575 837 579 841
rect 611 837 615 841
rect 619 837 623 841
rect 655 837 659 841
rect 663 837 667 841
rect 699 837 703 841
rect 707 837 711 841
rect 743 837 747 841
rect 751 837 755 841
rect 787 837 791 841
rect 795 837 799 841
rect 831 837 835 841
rect -367 810 -362 815
rect -348 810 -343 815
rect -336 810 -331 815
rect -317 810 -312 815
rect -303 810 -298 815
rect -284 810 -279 815
rect -351 524 -347 528
rect -328 524 -324 528
rect -317 524 -313 528
rect -294 524 -290 528
rect -284 524 -280 528
rect -261 524 -257 528
rect -252 524 -248 528
rect -229 524 -225 528
rect -220 524 -216 528
rect -197 524 -193 528
rect -188 524 -184 528
rect -165 524 -161 528
rect -352 277 -348 281
rect -329 277 -325 281
rect -318 277 -314 281
rect -295 277 -291 281
rect -285 277 -281 281
rect -262 277 -258 281
rect -253 277 -249 281
rect -230 277 -226 281
rect -221 277 -217 281
rect -198 277 -194 281
rect -189 277 -185 281
rect -166 277 -162 281
rect 2 217 6 221
rect 38 217 42 221
rect 46 217 50 221
rect 82 217 86 221
rect 90 217 94 221
rect 126 217 130 221
rect 134 217 138 221
rect 170 217 174 221
rect 178 217 182 221
rect 214 217 218 221
rect 222 217 226 221
rect 258 217 262 221
rect -348 51 -344 55
rect -325 51 -321 55
rect -314 51 -310 55
rect -291 51 -287 55
rect -281 51 -277 55
rect -258 51 -254 55
rect -249 51 -245 55
rect -226 51 -222 55
rect -217 51 -213 55
rect -194 51 -190 55
rect -185 51 -181 55
rect -162 51 -158 55
rect -351 -156 -347 -152
rect -328 -156 -324 -152
rect -317 -156 -313 -152
rect -294 -156 -290 -152
rect -284 -156 -280 -152
rect -261 -156 -257 -152
rect -252 -156 -248 -152
rect -229 -156 -225 -152
rect -220 -156 -216 -152
rect -197 -156 -193 -152
rect -188 -156 -184 -152
rect -165 -156 -161 -152
<< pdcontact >>
rect -331 1137 -327 1141
rect -283 1137 -279 1141
rect 194 1138 198 1142
rect -61 1132 -57 1136
rect -13 1132 -9 1136
rect 242 1138 246 1142
rect 462 1138 466 1142
rect 510 1138 514 1142
rect 1018 990 1022 994
rect 1043 990 1047 994
rect 1052 990 1056 994
rect 1077 990 1081 994
rect 1085 990 1089 994
rect 1110 990 1114 994
rect 1118 990 1122 994
rect 1143 990 1147 994
rect 1151 990 1155 994
rect 1176 990 1180 994
rect -189 940 -185 944
rect -153 940 -149 944
rect -145 940 -141 944
rect -109 940 -105 944
rect -101 940 -97 944
rect -65 940 -61 944
rect -57 940 -53 944
rect -21 940 -17 944
rect -13 940 -9 944
rect 23 940 27 944
rect 31 940 35 944
rect 67 940 71 944
rect 193 940 197 944
rect 229 940 233 944
rect 237 940 241 944
rect 273 940 277 944
rect 281 940 285 944
rect 317 940 321 944
rect 325 940 329 944
rect 361 940 365 944
rect 369 940 373 944
rect 405 940 409 944
rect 413 940 417 944
rect 449 940 453 944
rect 575 940 579 944
rect 611 940 615 944
rect 619 940 623 944
rect 655 940 659 944
rect 663 940 667 944
rect 699 940 703 944
rect 707 940 711 944
rect 743 940 747 944
rect 751 940 755 944
rect 787 940 791 944
rect 795 940 799 944
rect 831 940 835 944
rect -367 868 -362 873
rect -348 868 -343 873
rect -336 868 -331 873
rect -317 868 -312 873
rect -303 868 -298 873
rect -284 868 -279 873
rect -351 613 -347 617
rect -328 613 -324 617
rect -317 613 -313 617
rect -294 613 -290 617
rect -284 613 -280 617
rect -261 613 -257 617
rect -252 613 -248 617
rect -229 613 -225 617
rect -220 613 -216 617
rect -197 613 -193 617
rect -188 613 -184 617
rect -165 613 -161 617
rect -352 366 -348 370
rect -329 366 -325 370
rect -318 366 -314 370
rect -295 366 -291 370
rect -285 366 -281 370
rect -262 366 -258 370
rect -253 366 -249 370
rect -230 366 -226 370
rect -221 366 -217 370
rect -198 366 -194 370
rect -189 366 -185 370
rect -166 366 -162 370
rect 2 320 6 324
rect 38 320 42 324
rect 46 320 50 324
rect 82 320 86 324
rect 90 320 94 324
rect 126 320 130 324
rect 134 320 138 324
rect 170 320 174 324
rect 178 320 182 324
rect 214 320 218 324
rect 222 320 226 324
rect 258 320 262 324
rect -348 140 -344 144
rect -325 140 -321 144
rect -314 140 -310 144
rect -291 140 -287 144
rect -281 140 -277 144
rect -258 140 -254 144
rect -249 140 -245 144
rect -226 140 -222 144
rect -217 140 -213 144
rect -194 140 -190 144
rect -185 140 -181 144
rect -162 140 -158 144
rect -351 -67 -347 -63
rect -328 -67 -324 -63
rect -317 -67 -313 -63
rect -294 -67 -290 -63
rect -284 -67 -280 -63
rect -261 -67 -257 -63
rect -252 -67 -248 -63
rect -229 -67 -225 -63
rect -220 -67 -216 -63
rect -197 -67 -193 -63
rect -188 -67 -184 -63
rect -165 -67 -161 -63
<< polysilicon >>
rect -307 1141 -303 1153
rect -37 1136 -33 1148
rect 218 1142 222 1154
rect 486 1142 490 1154
rect -307 1103 -303 1131
rect -37 1098 -33 1126
rect 218 1104 222 1132
rect 486 1104 490 1132
rect -307 1074 -303 1089
rect -37 1069 -33 1084
rect 218 1075 222 1090
rect 486 1075 490 1090
rect 1030 994 1034 1004
rect 1065 994 1069 1004
rect 1098 994 1102 1004
rect 1131 994 1135 1004
rect 1164 994 1168 1004
rect -173 944 -169 949
rect -127 944 -123 949
rect -82 944 -78 949
rect -39 944 -35 949
rect 6 944 10 949
rect 49 944 53 949
rect 209 944 213 949
rect 255 944 259 949
rect 300 944 304 949
rect 343 944 347 949
rect 388 944 392 949
rect 431 944 435 949
rect 591 944 595 949
rect 637 944 641 949
rect 682 944 686 949
rect 725 944 729 949
rect 770 944 774 949
rect 813 944 817 949
rect -358 873 -354 879
rect -326 873 -322 877
rect -292 873 -288 877
rect -358 830 -354 864
rect -357 825 -354 830
rect -358 815 -354 825
rect -326 815 -322 864
rect -292 815 -288 864
rect -173 841 -169 933
rect -127 886 -123 933
rect -128 877 -123 886
rect -82 885 -78 933
rect -39 885 -35 933
rect -127 841 -123 877
rect -80 876 -78 885
rect -37 876 -35 885
rect 6 883 10 933
rect -82 841 -78 876
rect -39 841 -35 876
rect 7 874 10 883
rect 6 841 10 874
rect 49 841 53 933
rect 209 841 213 933
rect 255 886 259 933
rect 254 877 259 886
rect 300 885 304 933
rect 343 885 347 933
rect 255 841 259 877
rect 302 876 304 885
rect 345 876 347 885
rect 388 883 392 933
rect 300 841 304 876
rect 343 841 347 876
rect 389 874 392 883
rect 388 841 392 874
rect 431 841 435 933
rect 591 841 595 933
rect 637 886 641 933
rect 636 877 641 886
rect 682 885 686 933
rect 725 885 729 933
rect 637 841 641 877
rect 684 876 686 885
rect 727 876 729 885
rect 770 883 774 933
rect 682 841 686 876
rect 725 841 729 876
rect 771 874 774 883
rect 770 841 774 874
rect 813 841 817 933
rect 1030 912 1034 985
rect 1065 912 1069 985
rect 1098 912 1102 985
rect 1131 912 1135 985
rect 1164 912 1168 985
rect 1030 899 1034 903
rect 1065 899 1069 903
rect 1098 899 1102 903
rect 1131 899 1135 903
rect 1164 899 1168 903
rect -173 823 -169 830
rect -127 823 -123 830
rect -82 823 -78 830
rect -39 823 -35 830
rect 6 823 10 830
rect 49 823 53 830
rect 209 823 213 830
rect 255 823 259 830
rect 300 823 304 830
rect 343 823 347 830
rect 388 823 392 830
rect 431 823 435 830
rect 591 823 595 830
rect 637 823 641 830
rect 682 823 686 830
rect 725 823 729 830
rect 770 823 774 830
rect 813 823 817 830
rect -358 803 -354 806
rect -326 803 -322 806
rect -292 803 -288 806
rect -306 643 -205 646
rect -341 617 -338 626
rect -306 617 -303 643
rect -271 617 -268 626
rect -239 617 -236 626
rect -208 617 -205 643
rect -175 617 -172 626
rect -341 528 -338 611
rect -306 528 -303 611
rect -271 528 -268 611
rect -239 528 -236 611
rect -208 528 -205 611
rect -175 528 -172 611
rect -341 511 -338 522
rect -306 514 -303 522
rect -271 511 -268 522
rect -239 514 -236 522
rect -208 514 -205 522
rect -175 514 -172 522
rect -341 509 -268 511
rect -307 396 -206 399
rect -342 370 -339 379
rect -307 370 -304 396
rect -272 370 -269 379
rect -240 370 -237 379
rect -209 370 -206 396
rect -176 370 -173 379
rect -342 281 -339 364
rect -307 281 -304 364
rect -272 281 -269 364
rect -240 281 -237 364
rect -209 281 -206 364
rect -176 281 -173 364
rect 18 324 22 329
rect 64 324 68 329
rect 109 324 113 329
rect 152 324 156 329
rect 197 324 201 329
rect 240 324 244 329
rect -342 264 -339 275
rect -307 267 -304 275
rect -272 264 -269 275
rect -240 267 -237 275
rect -209 267 -206 275
rect -176 267 -173 275
rect -342 262 -269 264
rect 18 221 22 313
rect 64 266 68 313
rect 63 257 68 266
rect 109 265 113 313
rect 152 265 156 313
rect 64 221 68 257
rect 111 256 113 265
rect 154 256 156 265
rect 197 263 201 313
rect 109 221 113 256
rect 152 221 156 256
rect 198 254 201 263
rect 197 221 201 254
rect 240 221 244 313
rect 18 203 22 210
rect 64 203 68 210
rect 109 203 113 210
rect 152 203 156 210
rect 197 203 201 210
rect 240 203 244 210
rect -303 170 -202 173
rect -338 144 -335 153
rect -303 144 -300 170
rect -268 144 -265 153
rect -236 144 -233 153
rect -205 144 -202 170
rect -172 144 -169 153
rect -338 55 -335 138
rect -303 55 -300 138
rect -268 55 -265 138
rect -236 55 -233 138
rect -205 55 -202 138
rect -172 55 -169 138
rect -338 38 -335 49
rect -303 41 -300 49
rect -268 38 -265 49
rect -236 41 -233 49
rect -205 41 -202 49
rect -172 41 -169 49
rect -338 36 -265 38
rect -306 -37 -205 -34
rect -341 -63 -338 -54
rect -306 -63 -303 -37
rect -271 -63 -268 -54
rect -239 -63 -236 -54
rect -208 -63 -205 -37
rect -175 -63 -172 -54
rect -341 -152 -338 -69
rect -306 -152 -303 -69
rect -271 -152 -268 -69
rect -239 -152 -236 -69
rect -208 -152 -205 -69
rect -175 -152 -172 -69
rect -341 -169 -338 -158
rect -306 -166 -303 -158
rect -271 -169 -268 -158
rect -239 -166 -236 -158
rect -208 -166 -205 -158
rect -175 -166 -172 -158
rect -341 -171 -268 -169
<< polycontact >>
rect -313 1116 -307 1120
rect -43 1111 -37 1115
rect 212 1117 218 1121
rect 480 1117 486 1121
rect 1026 946 1030 950
rect -182 878 -173 887
rect -361 825 -357 830
rect -330 825 -326 830
rect -298 838 -292 844
rect -137 877 -128 886
rect -89 876 -80 885
rect -46 876 -37 885
rect -2 874 7 883
rect 39 882 49 891
rect 200 878 209 887
rect 245 877 254 886
rect 293 876 302 885
rect 336 876 345 885
rect 380 874 389 883
rect 421 882 431 891
rect 582 878 591 887
rect 627 877 636 886
rect 675 876 684 885
rect 718 876 727 885
rect 762 874 771 883
rect 803 882 813 891
rect 1061 945 1065 949
rect 1094 944 1098 948
rect 1127 943 1131 947
rect 1159 945 1164 949
rect -348 573 -341 579
rect -312 572 -306 578
rect -245 572 -239 578
rect -181 548 -175 553
rect -349 326 -342 332
rect -313 325 -307 331
rect -246 325 -240 331
rect -182 301 -176 306
rect 9 258 18 267
rect 54 257 63 266
rect 102 256 111 265
rect 145 256 154 265
rect 189 254 198 263
rect 230 262 240 271
rect -345 100 -338 106
rect -309 99 -303 105
rect -242 99 -236 105
rect -178 75 -172 80
rect -348 -107 -341 -101
rect -312 -108 -306 -102
rect -245 -108 -239 -102
rect -181 -132 -175 -127
<< metal1 >>
rect -392 1179 -234 1185
rect -392 831 -385 1179
rect -349 1162 -253 1163
rect -349 1161 -263 1162
rect -375 1154 -263 1161
rect -375 968 -366 1154
rect -349 1153 -253 1154
rect -331 1141 -327 1153
rect -318 1116 -313 1120
rect -283 1119 -279 1137
rect -238 1119 -234 1179
rect 176 1161 272 1164
rect 444 1161 540 1164
rect 176 1159 540 1161
rect 11 1158 540 1159
rect -71 1156 540 1158
rect -71 1155 272 1156
rect -71 1150 17 1155
rect 176 1154 272 1155
rect 444 1154 540 1156
rect -79 1148 17 1150
rect -61 1136 -57 1148
rect 194 1142 198 1154
rect 462 1142 466 1154
rect -283 1113 -234 1119
rect -283 1103 -279 1113
rect -48 1111 -43 1115
rect -13 1114 -9 1132
rect 207 1117 212 1121
rect 242 1120 246 1138
rect 242 1114 290 1120
rect 475 1117 480 1121
rect 510 1120 514 1138
rect -13 1108 -10 1114
rect -331 1074 -327 1099
rect -13 1098 -9 1108
rect 242 1104 246 1114
rect 510 1113 513 1120
rect 510 1104 514 1113
rect -350 1069 -272 1074
rect -260 1069 -253 1074
rect -61 1069 -57 1094
rect 194 1075 198 1100
rect 462 1075 466 1100
rect 175 1071 540 1075
rect 175 1070 272 1071
rect 14 1069 272 1070
rect 443 1069 540 1071
rect -350 1068 -253 1069
rect -80 1068 197 1069
rect -257 1066 197 1068
rect -257 1064 17 1066
rect -80 1063 17 1064
rect 821 1065 827 1072
rect 821 1060 1019 1065
rect 821 971 827 1060
rect 1015 1017 1020 1060
rect 1006 1009 1192 1017
rect 1018 994 1022 1009
rect 1151 994 1155 1009
rect 1047 990 1052 994
rect 1081 990 1085 994
rect 1114 990 1118 994
rect -196 970 94 971
rect -196 969 96 970
rect 186 969 844 971
rect -196 968 844 969
rect -375 966 844 968
rect -375 964 475 966
rect -375 963 96 964
rect -375 889 -366 963
rect -196 957 96 963
rect -196 956 80 957
rect -189 944 -185 956
rect -145 944 -141 956
rect -101 944 -97 956
rect -57 944 -53 956
rect -13 944 -9 956
rect 31 944 35 956
rect -153 929 -149 940
rect -109 929 -105 940
rect -65 929 -61 940
rect -21 929 -17 940
rect 23 929 27 940
rect -153 925 27 929
rect 23 891 32 925
rect 67 894 71 940
rect 86 912 96 957
rect 186 957 475 964
rect 482 963 844 966
rect 482 957 483 963
rect 186 956 462 957
rect 568 956 844 963
rect 193 944 197 956
rect 237 944 241 956
rect 281 944 285 956
rect 325 944 329 956
rect 369 944 373 956
rect 413 944 417 956
rect 575 944 579 956
rect 619 944 623 956
rect 663 944 667 956
rect 707 944 711 956
rect 751 944 755 956
rect 795 944 799 956
rect 997 949 1003 950
rect 1022 949 1026 950
rect 997 944 1026 949
rect 1059 945 1061 949
rect 229 929 233 940
rect 273 929 277 940
rect 317 929 321 940
rect 361 929 365 940
rect 405 929 409 940
rect 229 925 409 929
rect 67 893 79 894
rect -375 882 -271 889
rect -367 873 -362 882
rect -336 873 -331 882
rect -303 873 -298 882
rect -194 878 -182 887
rect -146 877 -137 886
rect -98 876 -89 885
rect -52 876 -46 885
rect -5 874 -2 883
rect 23 882 39 891
rect -348 844 -343 868
rect -317 844 -312 868
rect -348 838 -298 844
rect -284 841 -279 868
rect 23 841 27 882
rect 67 841 71 893
rect 78 882 79 893
rect 405 891 414 925
rect 449 894 453 940
rect 611 929 615 940
rect 655 929 659 940
rect 699 929 703 940
rect 743 929 747 940
rect 787 929 791 940
rect 611 925 791 929
rect 449 893 461 894
rect 191 885 200 887
rect 196 879 200 885
rect 191 878 200 879
rect 236 884 245 886
rect 241 878 245 884
rect 236 877 245 878
rect 287 876 293 885
rect 327 876 336 885
rect 371 882 380 883
rect 375 875 380 882
rect 371 874 380 875
rect 405 882 421 891
rect 449 882 456 893
rect 787 891 796 925
rect 831 894 835 940
rect 831 893 843 894
rect 405 841 409 882
rect 449 841 453 882
rect 579 878 582 887
rect 623 877 627 886
rect 672 876 675 885
rect 715 876 718 885
rect 753 874 762 883
rect 787 882 803 891
rect 831 883 837 893
rect 831 882 843 883
rect 787 841 791 882
rect 831 841 835 882
rect -392 830 -366 831
rect -392 825 -361 830
rect -336 829 -330 830
rect -338 825 -330 829
rect -317 815 -312 838
rect -284 835 -242 841
rect -149 837 -145 841
rect -105 837 -101 841
rect -61 837 -57 841
rect -17 837 -13 841
rect 233 837 237 841
rect 277 837 281 841
rect 321 837 325 841
rect 365 837 369 841
rect 615 837 619 841
rect 659 837 663 841
rect 703 837 707 841
rect 747 837 751 841
rect -284 815 -279 835
rect -343 810 -336 815
rect -367 806 -362 810
rect -303 806 -298 810
rect -373 805 -271 806
rect -365 799 -271 805
rect -246 741 -243 835
rect -232 818 -231 821
rect -189 823 -185 837
rect 31 823 35 837
rect 193 823 197 837
rect 413 823 417 837
rect 575 823 579 837
rect 795 823 799 837
rect -192 821 84 823
rect -226 818 84 821
rect -192 812 84 818
rect 190 814 466 823
rect 572 814 848 823
rect 190 812 848 814
rect -192 810 848 812
rect -192 808 466 810
rect 572 808 848 810
rect 997 741 1003 944
rect 1143 949 1147 990
rect 1176 949 1180 990
rect 1090 948 1093 949
rect 1090 944 1094 948
rect 1090 943 1093 944
rect 1125 943 1127 947
rect 1143 945 1159 949
rect 1176 945 1189 949
rect 1143 933 1147 945
rect 1043 929 1147 933
rect 1043 912 1047 929
rect 1077 912 1081 929
rect 1110 912 1114 929
rect 1143 912 1147 929
rect 1176 912 1180 945
rect 1018 900 1022 908
rect 1052 900 1056 908
rect 1085 900 1089 908
rect 1118 900 1122 908
rect 1151 900 1155 908
rect 1015 892 1201 900
rect -246 740 -216 741
rect -203 740 1003 741
rect -246 736 1003 740
rect -246 735 -216 736
rect -203 735 1003 736
rect -121 692 411 693
rect -198 687 411 692
rect -369 661 -205 662
rect -432 415 -425 661
rect -416 650 54 661
rect -351 617 -347 650
rect -317 617 -313 650
rect -284 617 -280 650
rect -252 617 -248 650
rect -229 649 54 650
rect -197 636 -133 642
rect -197 617 -193 636
rect -165 617 -161 636
rect -356 573 -348 579
rect -328 528 -324 613
rect -294 578 -290 613
rect -261 589 -257 613
rect -229 589 -225 613
rect -220 589 -216 613
rect -188 589 -184 613
rect -137 592 -133 636
rect -261 585 -184 589
rect -138 587 -21 592
rect -319 572 -312 578
rect -294 572 -245 578
rect -294 528 -290 572
rect -185 548 -181 553
rect -137 543 -133 587
rect -229 539 -133 543
rect -229 528 -225 539
rect -165 528 -161 539
rect -257 524 -252 528
rect -193 524 -188 528
rect -351 507 -347 524
rect -317 507 -313 524
rect -284 507 -280 524
rect -220 507 -216 524
rect -358 492 -201 507
rect -432 404 -206 415
rect -432 189 -425 404
rect -370 403 -206 404
rect -352 370 -348 403
rect -318 370 -314 403
rect -285 370 -281 403
rect -253 370 -249 403
rect -198 389 -133 395
rect -198 370 -194 389
rect -166 370 -162 389
rect -357 326 -349 332
rect -329 281 -325 366
rect -295 331 -291 366
rect -262 342 -258 366
rect -230 342 -226 366
rect -221 342 -217 366
rect -189 342 -185 366
rect -262 338 -185 342
rect -320 325 -313 331
rect -295 325 -246 331
rect -295 281 -291 325
rect -138 318 -133 389
rect -94 318 -83 463
rect -46 318 -39 319
rect -139 313 -39 318
rect -186 301 -182 306
rect -138 296 -133 313
rect -94 312 -83 313
rect -230 292 -133 296
rect -46 293 -39 313
rect -230 281 -226 292
rect -166 281 -162 292
rect -258 277 -253 281
rect -194 277 -189 281
rect -352 260 -348 277
rect -318 260 -314 277
rect -285 260 -281 277
rect -221 261 -217 277
rect -24 266 -21 587
rect 45 351 54 649
rect 397 612 409 687
rect 79 467 356 476
rect -5 342 297 351
rect -5 336 271 342
rect 2 324 6 336
rect 46 324 50 336
rect 90 324 94 336
rect 134 324 138 336
rect 178 324 182 336
rect 222 324 226 336
rect 38 309 42 320
rect 82 309 86 320
rect 126 309 130 320
rect 170 309 174 320
rect 214 309 218 320
rect 38 305 218 309
rect 214 271 223 305
rect 258 274 262 320
rect 289 296 296 342
rect 394 283 409 612
rect 712 283 727 673
rect 0 266 9 267
rect -222 260 -62 261
rect -352 245 -62 260
rect -24 258 9 266
rect 50 257 54 266
rect 99 256 102 265
rect 140 256 145 265
rect 184 255 189 263
rect 180 254 189 255
rect 214 262 230 271
rect 258 262 270 274
rect 394 271 731 283
rect -222 244 -62 245
rect -70 202 -62 244
rect 214 221 218 262
rect 258 221 262 262
rect 42 217 46 221
rect 86 217 90 221
rect 130 217 134 221
rect 174 217 178 221
rect 2 203 6 217
rect 222 203 226 217
rect -1 202 275 203
rect -432 178 -202 189
rect -70 188 275 202
rect -432 135 -425 178
rect -366 177 -202 178
rect -348 144 -344 177
rect -314 144 -310 177
rect -281 144 -277 177
rect -249 144 -245 177
rect -194 163 -129 169
rect -194 144 -190 163
rect -162 144 -158 163
rect -433 -18 -425 135
rect -353 100 -345 106
rect -325 55 -321 140
rect -291 105 -287 140
rect -258 116 -254 140
rect -226 116 -222 140
rect -134 160 -129 163
rect -134 154 90 160
rect -217 116 -213 140
rect -185 116 -181 140
rect -258 112 -181 116
rect -316 99 -309 105
rect -291 99 -242 105
rect -291 55 -287 99
rect -182 75 -178 80
rect -134 70 -129 154
rect -226 66 -129 70
rect -226 55 -222 66
rect -162 55 -158 66
rect -254 51 -249 55
rect -190 51 -185 55
rect -348 34 -344 51
rect -314 34 -310 51
rect -281 34 -277 51
rect -217 34 -213 51
rect -346 19 -198 34
rect 131 -14 143 153
rect 394 0 409 271
rect 712 270 727 271
rect 394 -14 408 0
rect -433 -29 -205 -18
rect -369 -30 -205 -29
rect -351 -63 -347 -30
rect -317 -63 -313 -30
rect -284 -63 -280 -30
rect -252 -63 -248 -30
rect 131 -31 408 -14
rect -197 -44 -131 -38
rect -197 -63 -193 -44
rect -165 -63 -161 -44
rect -356 -107 -348 -101
rect -328 -152 -324 -67
rect -294 -102 -290 -67
rect -261 -91 -257 -67
rect -229 -91 -225 -67
rect -220 -91 -216 -67
rect -188 -91 -184 -67
rect -261 -95 -184 -91
rect -137 -83 -132 -44
rect 131 -83 143 -31
rect 394 -32 408 -31
rect -137 -92 143 -83
rect -319 -108 -312 -102
rect -294 -108 -245 -102
rect -294 -152 -290 -108
rect -185 -132 -181 -127
rect -137 -137 -132 -92
rect -229 -141 -131 -137
rect -229 -152 -225 -141
rect -165 -152 -161 -141
rect -257 -156 -252 -152
rect -193 -156 -188 -152
rect -351 -172 -347 -156
rect -348 -173 -347 -172
rect -317 -173 -313 -156
rect -284 -173 -280 -156
rect -220 -173 -216 -156
rect -348 -179 -201 -173
rect 1125 -179 1130 892
rect -348 -188 1130 -179
rect -220 -189 1130 -188
rect -220 -191 1129 -189
<< m2contact >>
rect -263 1154 -253 1162
rect -81 1150 -71 1158
rect 290 1114 296 1120
rect -10 1108 -1 1114
rect 513 1113 523 1120
rect -272 1069 -260 1076
rect 475 957 482 966
rect 1054 945 1059 952
rect 86 903 96 912
rect -207 876 -194 887
rect -158 877 -146 886
rect -62 876 -52 885
rect -15 874 -5 883
rect 71 882 78 893
rect 190 879 196 885
rect 234 878 241 884
rect 277 874 287 886
rect 366 875 375 882
rect 456 882 465 893
rect 567 878 579 887
rect 612 877 623 886
rect 661 876 672 887
rect 707 876 715 885
rect 837 883 848 893
rect -377 798 -365 805
rect -271 799 -259 806
rect -231 814 -226 829
rect 1084 942 1090 952
rect 1119 943 1125 949
rect 1111 880 1121 887
rect -211 685 -198 696
rect -425 650 -416 661
rect -324 548 -316 553
rect -192 548 -185 553
rect -379 491 -358 508
rect -95 463 -78 482
rect -325 301 -317 306
rect -193 301 -186 306
rect -46 277 -39 293
rect -371 245 -352 261
rect 66 467 79 478
rect 356 465 373 482
rect 289 282 297 296
rect 712 673 727 693
rect 38 257 50 267
rect 90 255 99 266
rect 131 255 140 265
rect 176 255 184 269
rect 90 154 100 168
rect -321 75 -313 80
rect -189 75 -182 80
rect 130 153 144 171
rect -365 18 -346 34
rect -324 -132 -316 -127
rect -192 -132 -185 -127
rect -367 -188 -348 -172
<< metal2 >>
rect -159 1219 -154 1239
rect -423 1217 -154 1219
rect -425 1206 -154 1217
rect -425 661 -418 1206
rect -159 1202 -154 1206
rect -160 1194 -154 1202
rect -160 1158 -155 1194
rect -253 1154 -81 1158
rect -1 1108 46 1113
rect -9 1107 46 1108
rect -267 821 -263 1069
rect 41 1022 46 1107
rect 293 1055 296 1114
rect 523 1114 555 1119
rect 164 1050 296 1055
rect -158 1016 46 1022
rect 128 1021 135 1023
rect -208 876 -207 881
rect -158 886 -153 1016
rect -13 911 -9 912
rect -58 907 86 911
rect -58 885 -54 907
rect -13 883 -9 907
rect -208 855 -201 876
rect 128 887 135 1008
rect 78 882 135 887
rect 71 881 135 882
rect 164 883 167 1050
rect 477 907 482 957
rect 366 900 482 907
rect 164 879 190 883
rect 234 855 237 878
rect -208 852 237 855
rect 366 882 370 900
rect 551 885 555 1114
rect 935 963 943 1008
rect 935 955 1058 963
rect 1054 952 1058 955
rect 465 882 503 885
rect 366 874 370 875
rect -267 818 -231 821
rect -391 805 -372 808
rect -267 806 -263 818
rect -391 798 -377 805
rect -391 797 -372 798
rect -391 508 -385 797
rect -208 696 -201 852
rect 277 775 285 874
rect 272 774 285 775
rect 91 770 285 774
rect 498 772 502 882
rect 551 881 567 885
rect 91 634 97 770
rect 498 769 580 772
rect -316 548 -192 553
rect -391 494 -379 508
rect -389 491 -379 494
rect -389 481 -368 491
rect -388 255 -381 481
rect -78 467 66 474
rect -78 466 79 467
rect 91 391 98 634
rect 612 475 621 877
rect 848 883 930 887
rect 1085 884 1089 942
rect 1119 887 1122 943
rect 846 882 930 883
rect 373 465 622 475
rect 663 391 670 876
rect 712 693 715 876
rect 923 847 929 882
rect 1066 881 1089 884
rect 923 841 1021 847
rect 1066 776 1072 881
rect 1121 884 1122 887
rect 1111 848 1117 880
rect 91 382 677 391
rect -317 301 -193 306
rect -39 277 45 282
rect -46 276 45 277
rect 38 267 45 276
rect -388 246 -371 255
rect -388 32 -381 246
rect 91 266 98 382
rect 663 380 670 382
rect 176 282 289 289
rect 176 278 297 282
rect 176 269 184 278
rect 90 168 97 255
rect 134 171 138 255
rect -313 75 -189 80
rect -388 27 -376 32
rect -388 18 -365 27
rect -388 -180 -381 18
rect -316 -132 -192 -127
rect -388 -188 -367 -180
rect -388 -189 -363 -188
<< m3contact >>
rect 128 1008 138 1021
rect 933 1008 944 1017
rect 580 769 588 776
rect 1021 841 1032 851
rect 1111 841 1121 848
rect 1066 769 1072 776
<< metal3 >>
rect 138 1008 933 1017
rect 1032 841 1111 847
rect 588 769 1066 774
<< labels >>
rlabel metal1 261 268 261 268 1 node_c2
rlabel metal1 -279 495 -279 495 1 gnd
rlabel metal1 -364 654 -364 654 1 vdd
rlabel metal1 -316 -105 -316 -105 1 node_b3
rlabel metal1 -354 -104 -354 -104 1 node_a3
rlabel metal1 -312 101 -312 101 1 node_b2
rlabel metal1 -349 102 -349 102 1 node_a2
rlabel metal1 -318 328 -318 328 1 node_b1
rlabel metal1 -354 329 -354 329 1 node_a1
rlabel metal1 -316 576 -316 576 1 node_b0
rlabel metal1 -354 574 -354 574 1 node_a0
rlabel metal1 -148 838 -148 838 1 node_x
rlabel metal1 234 838 234 838 1 node_x
rlabel metal1 616 838 616 838 1 node_x
rlabel metal1 -316 1117 -316 1117 1 node_b3
rlabel metal1 -46 1113 -46 1113 1 node_b2
rlabel metal1 209 1119 209 1119 1 node_b1
rlabel metal1 476 1118 476 1118 1 node_b0
rlabel metal1 -335 828 -335 828 1 node_a3
rlabel metal1 -95 882 -95 882 1 node_a2
rlabel metal1 331 880 331 880 1 node_a1
rlabel metal1 757 875 757 875 1 node_a0
rlabel metal1 1183 947 1183 947 1 node_c1
<< end >>
