magic
tech scmos
timestamp 1700163268
<< nwell >>
rect -4 165 96 195
rect -195 141 -120 163
rect -2 64 98 94
rect 1 -35 101 -5
rect -197 -78 -122 -56
rect 3 -143 103 -113
<< ntransistor >>
rect 11 119 15 128
rect 43 119 47 128
rect 77 119 81 128
rect -161 105 -157 119
rect 13 18 17 27
rect 45 18 49 27
rect 79 18 83 27
rect 16 -81 20 -72
rect 48 -81 52 -72
rect 82 -81 86 -72
rect -163 -114 -159 -100
rect 18 -189 22 -180
rect 50 -189 54 -180
rect 84 -189 88 -180
<< ptransistor >>
rect 11 177 15 186
rect 43 177 47 186
rect 77 177 81 186
rect -161 147 -157 157
rect 13 76 17 85
rect 45 76 49 85
rect 79 76 83 85
rect 16 -23 20 -14
rect 48 -23 52 -14
rect 82 -23 86 -14
rect -163 -72 -159 -62
rect 18 -131 22 -122
rect 50 -131 54 -122
rect 84 -131 88 -122
<< ndiffusion >>
rect 7 123 11 128
rect 2 119 11 123
rect 15 123 21 128
rect 15 119 26 123
rect 38 123 43 128
rect 33 119 43 123
rect 47 123 52 128
rect 47 119 57 123
rect 71 123 77 128
rect 66 119 77 123
rect 81 123 85 128
rect 81 119 90 123
rect -181 115 -161 119
rect -185 105 -161 115
rect -157 115 -137 119
rect -157 105 -133 115
rect 9 22 13 27
rect 4 18 13 22
rect 17 22 23 27
rect 17 18 28 22
rect 40 22 45 27
rect 35 18 45 22
rect 49 22 54 27
rect 49 18 59 22
rect 73 22 79 27
rect 68 18 79 22
rect 83 22 87 27
rect 83 18 92 22
rect 12 -77 16 -72
rect 7 -81 16 -77
rect 20 -77 26 -72
rect 20 -81 31 -77
rect 43 -77 48 -72
rect 38 -81 48 -77
rect 52 -77 57 -72
rect 52 -81 62 -77
rect 76 -77 82 -72
rect 71 -81 82 -77
rect 86 -77 90 -72
rect 86 -81 95 -77
rect -183 -104 -163 -100
rect -187 -114 -163 -104
rect -159 -104 -139 -100
rect -159 -114 -135 -104
rect 14 -185 18 -180
rect 9 -189 18 -185
rect 22 -185 28 -180
rect 22 -189 33 -185
rect 45 -185 50 -180
rect 40 -189 50 -185
rect 54 -185 59 -180
rect 54 -189 64 -185
rect 78 -185 84 -180
rect 73 -189 84 -185
rect 88 -185 92 -180
rect 88 -189 97 -185
<< pdiffusion >>
rect 7 181 11 186
rect 2 177 11 181
rect 15 181 21 186
rect 15 177 26 181
rect 38 181 43 186
rect 33 177 43 181
rect 47 181 52 186
rect 47 177 57 181
rect 71 181 77 186
rect 66 177 77 181
rect 81 181 85 186
rect 81 177 90 181
rect -181 153 -161 157
rect -185 147 -161 153
rect -157 153 -137 157
rect -157 147 -133 153
rect 9 80 13 85
rect 4 76 13 80
rect 17 80 23 85
rect 17 76 28 80
rect 40 80 45 85
rect 35 76 45 80
rect 49 80 54 85
rect 49 76 59 80
rect 73 80 79 85
rect 68 76 79 80
rect 83 80 87 85
rect 83 76 92 80
rect 12 -19 16 -14
rect 7 -23 16 -19
rect 20 -19 26 -14
rect 20 -23 31 -19
rect 43 -19 48 -14
rect 38 -23 48 -19
rect 52 -19 57 -14
rect 52 -23 62 -19
rect 76 -19 82 -14
rect 71 -23 82 -19
rect 86 -19 90 -14
rect 86 -23 95 -19
rect -183 -66 -163 -62
rect -187 -72 -163 -66
rect -159 -66 -139 -62
rect -159 -72 -135 -66
rect 14 -127 18 -122
rect 9 -131 18 -127
rect 22 -127 28 -122
rect 22 -131 33 -127
rect 45 -127 50 -122
rect 40 -131 50 -127
rect 54 -127 59 -122
rect 54 -131 64 -127
rect 78 -127 84 -122
rect 73 -131 84 -127
rect 88 -127 92 -122
rect 88 -131 97 -127
<< ndcontact >>
rect 2 123 7 128
rect 21 123 26 128
rect 33 123 38 128
rect 52 123 57 128
rect 66 123 71 128
rect 85 123 90 128
rect -185 115 -181 119
rect -137 115 -133 119
rect 4 22 9 27
rect 23 22 28 27
rect 35 22 40 27
rect 54 22 59 27
rect 68 22 73 27
rect 87 22 92 27
rect 7 -77 12 -72
rect 26 -77 31 -72
rect 38 -77 43 -72
rect 57 -77 62 -72
rect 71 -77 76 -72
rect 90 -77 95 -72
rect -187 -104 -183 -100
rect -139 -104 -135 -100
rect 9 -185 14 -180
rect 28 -185 33 -180
rect 40 -185 45 -180
rect 59 -185 64 -180
rect 73 -185 78 -180
rect 92 -185 97 -180
<< pdcontact >>
rect 2 181 7 186
rect 21 181 26 186
rect 33 181 38 186
rect 52 181 57 186
rect 66 181 71 186
rect 85 181 90 186
rect -185 153 -181 157
rect -137 153 -133 157
rect 4 80 9 85
rect 23 80 28 85
rect 35 80 40 85
rect 54 80 59 85
rect 68 80 73 85
rect 87 80 92 85
rect 7 -19 12 -14
rect 26 -19 31 -14
rect 38 -19 43 -14
rect 57 -19 62 -14
rect 71 -19 76 -14
rect 90 -19 95 -14
rect -187 -66 -183 -62
rect -139 -66 -135 -62
rect 9 -127 14 -122
rect 28 -127 33 -122
rect 40 -127 45 -122
rect 59 -127 64 -122
rect 73 -127 78 -122
rect 92 -127 97 -122
<< polysilicon >>
rect 11 186 15 192
rect 43 186 47 190
rect 77 186 81 190
rect -161 157 -157 169
rect -161 119 -157 147
rect 11 143 15 177
rect 12 138 15 143
rect 11 128 15 138
rect 43 128 47 177
rect 77 128 81 177
rect 11 116 15 119
rect 43 116 47 119
rect 77 116 81 119
rect -161 90 -157 105
rect 13 85 17 91
rect 45 85 49 89
rect 79 85 83 89
rect 13 42 17 76
rect 14 37 17 42
rect 13 27 17 37
rect 45 27 49 76
rect 79 27 83 76
rect 13 15 17 18
rect 45 15 49 18
rect 79 15 83 18
rect 16 -14 20 -8
rect 48 -14 52 -10
rect 82 -14 86 -10
rect -163 -62 -159 -50
rect 16 -57 20 -23
rect 17 -62 20 -57
rect 16 -72 20 -62
rect 48 -72 52 -23
rect 82 -72 86 -23
rect -163 -100 -159 -72
rect 16 -84 20 -81
rect 48 -84 52 -81
rect 82 -84 86 -81
rect -163 -129 -159 -114
rect 18 -122 22 -116
rect 50 -122 54 -118
rect 84 -122 88 -118
rect 18 -165 22 -131
rect 19 -170 22 -165
rect 18 -180 22 -170
rect 50 -180 54 -131
rect 84 -180 88 -131
rect 18 -192 22 -189
rect 50 -192 54 -189
rect 84 -192 88 -189
<< polycontact >>
rect -167 132 -161 136
rect 8 138 12 143
rect 39 138 43 143
rect 71 151 77 157
rect 10 37 14 42
rect 41 37 45 42
rect 73 50 79 56
rect 13 -62 17 -57
rect 44 -62 48 -57
rect 76 -49 82 -43
rect -169 -87 -163 -83
rect 15 -170 19 -165
rect 46 -170 50 -165
rect 78 -157 84 -151
<< metal1 >>
rect -42 195 133 201
rect -42 179 -33 195
rect 2 186 7 195
rect 33 186 38 195
rect 66 186 71 195
rect -257 169 -33 179
rect -257 167 -192 169
rect -257 -39 -250 167
rect -185 157 -181 169
rect 21 157 26 181
rect 52 157 57 181
rect -137 138 -133 153
rect 21 151 71 157
rect 85 154 90 181
rect 85 153 93 154
rect -47 138 8 143
rect 30 138 39 143
rect -220 132 -167 136
rect -137 134 -42 138
rect 30 137 43 138
rect 30 135 34 137
rect -220 29 -217 132
rect -137 119 -133 134
rect -185 90 -181 115
rect -204 82 -117 90
rect -107 82 -106 90
rect -204 80 -106 82
rect -95 29 -90 47
rect -220 26 -90 29
rect -257 -40 -195 -39
rect -257 -50 -107 -40
rect -86 -41 -83 134
rect -27 131 34 135
rect -27 97 -22 131
rect 52 128 57 151
rect 84 149 93 153
rect 85 128 90 149
rect 26 123 33 128
rect 2 119 7 123
rect 66 119 71 123
rect -4 112 93 119
rect 125 100 133 195
rect -62 92 -22 97
rect -3 94 133 100
rect -62 42 -57 92
rect 4 85 9 94
rect 35 85 40 94
rect 68 85 73 94
rect 23 56 28 80
rect 54 56 59 80
rect 23 50 73 56
rect 87 53 92 80
rect 87 52 95 53
rect -62 37 10 42
rect -187 -62 -183 -50
rect -224 -87 -169 -83
rect -139 -84 -135 -66
rect -62 -84 -57 37
rect 37 37 41 42
rect 37 36 45 37
rect 54 27 59 50
rect 86 48 95 52
rect 87 27 92 48
rect 28 22 35 27
rect 4 18 9 22
rect 68 18 73 22
rect -2 11 96 18
rect 125 1 133 94
rect 0 -5 133 1
rect 7 -14 12 -5
rect 38 -14 43 -5
rect 71 -14 76 -5
rect 26 -43 31 -19
rect 57 -43 62 -19
rect -42 -50 0 -47
rect 26 -49 76 -43
rect 90 -46 95 -19
rect 90 -47 98 -46
rect -3 -57 0 -50
rect -3 -62 13 -57
rect 57 -72 62 -49
rect 89 -51 98 -47
rect 90 -72 95 -51
rect 31 -77 38 -72
rect 7 -81 12 -77
rect 71 -81 76 -77
rect -224 -156 -220 -87
rect -139 -90 -57 -84
rect 1 -88 99 -81
rect -139 -100 -135 -90
rect -62 -100 41 -97
rect -187 -129 -183 -104
rect -206 -130 -108 -129
rect -206 -139 -120 -130
rect -109 -139 -108 -130
rect -62 -156 -57 -100
rect 125 -107 133 -5
rect 2 -113 133 -107
rect 9 -122 14 -113
rect 40 -122 45 -113
rect 73 -122 78 -113
rect -224 -161 -57 -156
rect 28 -151 33 -127
rect 59 -151 64 -127
rect 28 -157 78 -151
rect 92 -154 97 -127
rect 92 -155 100 -154
rect 11 -170 15 -165
rect 46 -165 50 -164
rect 46 -171 50 -170
rect 59 -180 64 -157
rect 91 -159 100 -155
rect 92 -180 97 -159
rect 33 -185 40 -180
rect 9 -189 14 -185
rect 73 -189 78 -185
rect 3 -196 101 -189
<< m2contact >>
rect -117 82 -107 90
rect -95 47 -90 55
rect 93 111 105 120
rect -86 -50 -78 -41
rect 28 36 37 42
rect 96 10 108 19
rect -50 -50 -42 -42
rect 99 -89 111 -80
rect 41 -100 47 -94
rect -120 -139 -109 -130
rect -1 -170 11 -165
rect 41 -171 46 -164
rect -8 -198 3 -189
rect 101 -197 113 -188
<< metal2 >>
rect 105 111 189 119
rect -115 -130 -110 82
rect -90 47 21 55
rect -78 -50 -50 -47
rect -114 -190 -109 -139
rect -37 -165 -34 47
rect 18 42 21 47
rect 18 36 28 42
rect 181 19 189 111
rect 108 11 189 19
rect 44 -94 47 -66
rect 181 -81 189 11
rect 111 -89 189 -81
rect 41 -164 44 -100
rect -37 -170 -1 -165
rect 181 -185 189 -89
rect 104 -188 190 -185
rect -114 -197 -8 -190
rect 113 -193 190 -188
<< labels >>
rlabel metal1 -90 174 -90 174 1 vdd
rlabel metal1 -131 -135 -131 -135 1 gnd
rlabel metal1 -187 134 -187 134 1 node_s0
rlabel metal1 -190 -86 -190 -86 1 node_s1
rlabel metal1 89 150 89 150 1 node_d0
rlabel metal1 90 50 90 50 1 node_d1
rlabel metal1 95 -49 95 -49 1 node_d2
rlabel metal1 97 -157 97 -157 1 node_d3
<< end >>
