magic
tech scmos
timestamp 1699126766
<< nwell >>
rect -735 299 -557 334
<< ntransistor >>
rect -716 231 -712 240
rect -681 231 -677 240
rect -648 231 -644 240
rect -615 231 -611 240
rect -582 231 -578 240
<< ptransistor >>
rect -716 313 -712 322
rect -681 313 -677 322
rect -648 313 -644 322
rect -615 313 -611 322
rect -582 313 -578 322
<< ndiffusion >>
rect -724 236 -716 240
rect -728 231 -716 236
rect -712 236 -703 240
rect -712 231 -699 236
rect -690 236 -681 240
rect -694 231 -681 236
rect -677 236 -669 240
rect -677 231 -665 236
rect -657 236 -648 240
rect -661 231 -648 236
rect -644 236 -636 240
rect -644 231 -632 236
rect -624 236 -615 240
rect -628 231 -615 236
rect -611 236 -603 240
rect -611 231 -599 236
rect -591 236 -582 240
rect -595 231 -582 236
rect -578 236 -570 240
rect -578 231 -566 236
<< pdiffusion >>
rect -724 318 -716 322
rect -728 313 -716 318
rect -712 318 -703 322
rect -712 313 -699 318
rect -690 318 -681 322
rect -694 313 -681 318
rect -677 318 -669 322
rect -677 313 -665 318
rect -657 318 -648 322
rect -661 313 -648 318
rect -644 318 -636 322
rect -644 313 -632 318
rect -624 318 -615 322
rect -628 313 -615 318
rect -611 318 -603 322
rect -611 313 -599 318
rect -591 318 -582 322
rect -595 313 -582 318
rect -578 318 -570 322
rect -578 313 -566 318
<< ndcontact >>
rect -728 236 -724 240
rect -703 236 -699 240
rect -694 236 -690 240
rect -669 236 -665 240
rect -661 236 -657 240
rect -636 236 -632 240
rect -628 236 -624 240
rect -603 236 -599 240
rect -595 236 -591 240
rect -570 236 -566 240
<< pdcontact >>
rect -728 318 -724 322
rect -703 318 -699 322
rect -694 318 -690 322
rect -669 318 -665 322
rect -661 318 -657 322
rect -636 318 -632 322
rect -628 318 -624 322
rect -603 318 -599 322
rect -595 318 -591 322
rect -570 318 -566 322
<< polysilicon >>
rect -716 322 -712 332
rect -681 322 -677 332
rect -648 322 -644 332
rect -615 322 -611 332
rect -582 322 -578 332
rect -716 240 -712 313
rect -681 240 -677 313
rect -648 240 -644 313
rect -615 240 -611 313
rect -582 240 -578 313
rect -716 227 -712 231
rect -681 227 -677 231
rect -648 227 -644 231
rect -615 227 -611 231
rect -582 227 -578 231
<< polycontact >>
rect -720 274 -716 278
rect -685 273 -681 277
rect -652 272 -648 276
rect -619 271 -615 275
rect -587 273 -582 277
<< metal1 >>
rect -740 337 -554 345
rect -728 322 -724 337
rect -595 322 -591 337
rect -699 318 -694 322
rect -665 318 -661 322
rect -632 318 -628 322
rect -724 274 -720 278
rect -603 277 -599 318
rect -570 277 -566 318
rect -689 273 -685 277
rect -656 272 -652 276
rect -623 271 -619 275
rect -603 273 -587 277
rect -570 273 -557 277
rect -603 261 -599 273
rect -703 257 -599 261
rect -703 240 -699 257
rect -669 240 -665 257
rect -636 240 -632 257
rect -603 240 -599 257
rect -570 240 -566 273
rect -728 228 -724 236
rect -694 228 -690 236
rect -661 228 -657 236
rect -628 228 -624 236
rect -595 228 -591 236
rect -731 220 -545 228
<< labels >>
rlabel metal1 -678 340 -678 340 5 vdd
rlabel metal1 -697 320 -697 320 1 node_x
rlabel metal1 -663 319 -663 319 1 node_y
rlabel metal1 -630 319 -630 319 1 node_m
rlabel metal1 -601 275 -601 275 1 node_nor
rlabel metal1 -567 274 -567 274 1 node_out
rlabel metal1 -722 276 -722 276 1 node_a
rlabel metal1 -688 274 -688 274 1 node_b
rlabel metal1 -655 275 -655 275 1 node_c
rlabel metal1 -621 273 -621 273 1 node_d
rlabel metal1 -668 224 -668 224 1 gnd
<< end >>
