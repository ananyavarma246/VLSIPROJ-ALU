magic
tech scmos
timestamp 1699686448
<< nwell >>
rect -497 396 -397 426
<< ntransistor >>
rect -482 350 -478 359
rect -450 350 -446 359
rect -416 350 -412 359
<< ptransistor >>
rect -482 408 -478 417
rect -450 408 -446 417
rect -416 408 -412 417
<< ndiffusion >>
rect -486 354 -482 359
rect -491 350 -482 354
rect -478 354 -472 359
rect -478 350 -467 354
rect -455 354 -450 359
rect -460 350 -450 354
rect -446 354 -441 359
rect -446 350 -436 354
rect -422 354 -416 359
rect -427 350 -416 354
rect -412 354 -408 359
rect -412 350 -403 354
<< pdiffusion >>
rect -486 412 -482 417
rect -491 408 -482 412
rect -478 412 -472 417
rect -478 408 -467 412
rect -455 412 -450 417
rect -460 408 -450 412
rect -446 412 -441 417
rect -446 408 -436 412
rect -422 412 -416 417
rect -427 408 -416 412
rect -412 412 -408 417
rect -412 408 -403 412
<< ndcontact >>
rect -491 354 -486 359
rect -472 354 -467 359
rect -460 354 -455 359
rect -441 354 -436 359
rect -427 354 -422 359
rect -408 354 -403 359
<< pdcontact >>
rect -491 412 -486 417
rect -472 412 -467 417
rect -460 412 -455 417
rect -441 412 -436 417
rect -427 412 -422 417
rect -408 412 -403 417
<< polysilicon >>
rect -482 417 -478 423
rect -450 417 -446 421
rect -416 417 -412 421
rect -482 374 -478 408
rect -481 369 -478 374
rect -482 359 -478 369
rect -450 359 -446 408
rect -416 359 -412 408
rect -482 347 -478 350
rect -450 347 -446 350
rect -416 347 -412 350
<< polycontact >>
rect -485 369 -481 374
rect -454 369 -450 374
rect -422 382 -416 388
<< metal1 >>
rect -498 426 -395 433
rect -491 417 -486 426
rect -460 417 -455 426
rect -427 417 -422 426
rect -472 388 -467 412
rect -441 388 -436 412
rect -472 382 -422 388
rect -408 385 -403 412
rect -491 369 -485 374
rect -460 369 -454 374
rect -441 359 -436 382
rect -408 380 -400 385
rect -408 359 -403 380
rect -467 354 -460 359
rect -491 350 -486 354
rect -427 350 -422 354
rect -497 343 -390 350
<< labels >>
rlabel metal1 -433 427 -433 427 1 vdd
rlabel metal1 -489 372 -489 372 1 node_a
rlabel metal1 -458 372 -458 372 1 node_b
rlabel metal1 -467 345 -467 345 1 gnd
rlabel metal1 -462 357 -462 357 1 node_x
rlabel metal1 -436 384 -436 384 1 node_inter
rlabel metal1 -404 383 -404 383 1 node_out
<< end >>
