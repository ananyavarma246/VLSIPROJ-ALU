magic
tech scmos
timestamp 1699098528
<< nwell >>
rect -2797 924 -2593 956
<< ntransistor >>
rect -2781 849 -2778 855
rect -2746 849 -2743 855
rect -2711 849 -2708 855
rect -2679 849 -2676 855
rect -2648 849 -2645 855
rect -2615 849 -2612 855
<< ptransistor >>
rect -2781 938 -2778 944
rect -2746 938 -2743 944
rect -2711 938 -2708 944
rect -2679 938 -2676 944
rect -2648 938 -2645 944
rect -2615 938 -2612 944
<< ndiffusion >>
rect -2787 851 -2781 855
rect -2791 849 -2781 851
rect -2778 851 -2768 855
rect -2778 849 -2764 851
rect -2753 851 -2746 855
rect -2757 849 -2746 851
rect -2743 851 -2734 855
rect -2743 849 -2730 851
rect -2720 851 -2711 855
rect -2724 849 -2711 851
rect -2708 851 -2701 855
rect -2708 849 -2697 851
rect -2688 851 -2679 855
rect -2692 849 -2679 851
rect -2676 851 -2669 855
rect -2676 849 -2665 851
rect -2656 851 -2648 855
rect -2660 849 -2648 851
rect -2645 851 -2637 855
rect -2645 849 -2633 851
rect -2624 851 -2615 855
rect -2628 849 -2615 851
rect -2612 851 -2605 855
rect -2612 849 -2601 851
<< pdiffusion >>
rect -2787 940 -2781 944
rect -2791 938 -2781 940
rect -2778 940 -2768 944
rect -2778 938 -2764 940
rect -2753 940 -2746 944
rect -2757 938 -2746 940
rect -2743 940 -2734 944
rect -2743 938 -2730 940
rect -2720 940 -2711 944
rect -2724 938 -2711 940
rect -2708 940 -2701 944
rect -2708 938 -2697 940
rect -2688 940 -2679 944
rect -2692 938 -2679 940
rect -2676 940 -2669 944
rect -2676 938 -2665 940
rect -2656 940 -2648 944
rect -2660 938 -2648 940
rect -2645 940 -2637 944
rect -2645 938 -2633 940
rect -2624 940 -2615 944
rect -2628 938 -2615 940
rect -2612 940 -2605 944
rect -2612 938 -2601 940
<< ndcontact >>
rect -2791 851 -2787 855
rect -2768 851 -2764 855
rect -2757 851 -2753 855
rect -2734 851 -2730 855
rect -2724 851 -2720 855
rect -2701 851 -2697 855
rect -2692 851 -2688 855
rect -2669 851 -2665 855
rect -2660 851 -2656 855
rect -2637 851 -2633 855
rect -2628 851 -2624 855
rect -2605 851 -2601 855
<< pdcontact >>
rect -2791 940 -2787 944
rect -2768 940 -2764 944
rect -2757 940 -2753 944
rect -2734 940 -2730 944
rect -2724 940 -2720 944
rect -2701 940 -2697 944
rect -2692 940 -2688 944
rect -2669 940 -2665 944
rect -2660 940 -2656 944
rect -2637 940 -2633 944
rect -2628 940 -2624 944
rect -2605 940 -2601 944
<< polysilicon >>
rect -2746 970 -2645 973
rect -2781 944 -2778 953
rect -2746 944 -2743 970
rect -2711 944 -2708 953
rect -2679 944 -2676 953
rect -2648 944 -2645 970
rect -2615 944 -2612 953
rect -2781 855 -2778 938
rect -2746 855 -2743 938
rect -2711 855 -2708 938
rect -2679 855 -2676 938
rect -2648 855 -2645 938
rect -2615 855 -2612 938
rect -2781 838 -2778 849
rect -2746 841 -2743 849
rect -2711 838 -2708 849
rect -2679 841 -2676 849
rect -2648 841 -2645 849
rect -2615 841 -2612 849
rect -2781 836 -2708 838
<< polycontact >>
rect -2788 900 -2781 906
rect -2752 899 -2746 905
rect -2685 899 -2679 905
rect -2621 875 -2615 880
<< metal1 >>
rect -2809 977 -2645 989
rect -2791 944 -2787 977
rect -2757 944 -2753 977
rect -2724 944 -2720 977
rect -2692 944 -2688 977
rect -2637 963 -2559 969
rect -2637 944 -2633 963
rect -2605 944 -2601 963
rect -2795 900 -2788 906
rect -2768 855 -2764 940
rect -2734 905 -2730 940
rect -2701 916 -2697 940
rect -2669 916 -2665 940
rect -2660 916 -2656 940
rect -2628 916 -2624 940
rect -2701 912 -2624 916
rect -2757 899 -2752 905
rect -2734 899 -2685 905
rect -2734 855 -2730 899
rect -2625 875 -2621 880
rect -2577 870 -2572 963
rect -2669 866 -2562 870
rect -2669 855 -2665 866
rect -2605 855 -2601 866
rect -2697 851 -2692 855
rect -2633 851 -2628 855
rect -2791 834 -2787 851
rect -2757 834 -2753 851
rect -2724 834 -2720 851
rect -2660 834 -2656 851
rect -2806 819 -2641 834
<< m2contact >>
rect -2764 875 -2756 880
rect -2632 875 -2625 880
<< metal2 >>
rect -2756 875 -2632 880
<< labels >>
rlabel metal1 -2715 985 -2715 985 5 vdd
rlabel metal1 -2792 903 -2792 903 1 node_a
rlabel metal1 -2755 902 -2755 902 1 node_b
rlabel metal1 -2766 902 -2766 902 1 node_anot
rlabel metal1 -2730 901 -2730 901 1 node_bnot
rlabel metal1 -2775 829 -2775 829 1 gnd
rlabel metal1 -2573 918 -2573 918 1 node_out
rlabel metal1 -2695 853 -2695 853 1 node_x
rlabel metal1 -2630 853 -2630 853 1 node_y
rlabel metal1 -2668 914 -2668 914 1 node_z
<< end >>
