.include TSMC_180nm.txt
.include addsub.sub



.param SUPPLY = 1.8
.param LAMBDA = 0.18u


.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param wn3 = {10*LAMBDA}
.param wn4 = {10*LAMBDA}
.param wn5 = {10*LAMBDA}
.param wn6 = {10*LAMBDA}
.param wn7 = {10*LAMBDA}

.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}
.param ln3 = {2*LAMBDA}
.param ln4 = {2*LAMBDA}
.param ln5 = {2*LAMBDA}
.param ln6 = {2*LAMBDA}
.param ln7 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param wp3 = wn1
.param wp4 = wn1
.param wp5 = wn1
.param wp6 = wn1
.param wp7 = wn1 

.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}
.param lp3 = {LAMBDA}
.param lp4 = {LAMBDA}
.param lp5 = {LAMBDA}
.param lp6 = {LAMBDA}
.param lp7 = {LAMBDA}

.global gnd

Vdd node_x gnd 'SUPPLY'

V_in_a0 node_a0 gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 50ns)
V_in_a1 node_a1 gnd PULSE(0 1.8 0ns 100ps 100ps 30ns 60ns)
V_in_a2 node_a2 gnd PULSE(0 1.8 0ns 100ps 100ps 40ns 70ns)
V_in_a3 node_a3 gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 80ns)

V_in_b0 node_b0 gnd PULSE(0 1.8 0ns 100ps 100ps 30ns 60ns)
V_in_b1 node_b1 gnd PULSE(0 1.8 0ns 100ps 100ps 40ns 70ns)
V_in_b2 node_b2 gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 80ns)
V_in_b3 node_b3 gnd PULSE(0 1.8 0ns 100ps 100ps 60ns 90ns)


V_in_c node_cin gnd PULSE(0 1.8 0ns 100ps 100ps 30ns 60ns)

X1 node_a0 node_a1 node_a2 node_a3 node_b0 node_b1 node_b2 node_b3 node_cin node_s1 node_s2 node_s3 node_s4 node_cout node_x gnd addsub


C1 node_s1 gnd 100f
C2 node_s2 gnd 100f
C3 node_s3 gnd 100f
C4 node_s4 gnd 100f
C5 node_cout gnd 100f

.tran 1n 800n

.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(node_a0) v(node_a1)+2  v(node_a2)+4 v(node_a3)+6 v(node_b0)+8 v(node_b1)+10  v(node_b2)+12 v(node_b3)+14 v(node_cin)+16 v(node_s1)+18 v(node_s2)+20 v(node_s3)+22 v(node_s4)+24 v(node_cout)+26
hardcopy image.ps v(node_a0) v(node_a1)+2  v(node_a2)+4 v(node_a3)+6 v(node_b0)+8 v(node_b1)+10  v(node_b2)+12 v(node_b3)+14 v(node_cin)+16 v(node_s1)+18 v(node_s2)+20 v(node_s3)+22 v(node_s4)+24 v(node_cout)+26
.end
.endc