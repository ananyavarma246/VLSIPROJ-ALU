//alu implementation
.include TSMC_180nm.txt

// including seperating blocks 

.include alu.sub


// parameters
.param SUPPLY = 1.8
.param LAMBDA = 0.18u


.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param wn3 = {10*LAMBDA}
.param wn4 = {10*LAMBDA}
.param wn5 = {10*LAMBDA}
.param wn6 = {10*LAMBDA}
.param wn7 = {10*LAMBDA}

.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}
.param ln3 = {2*LAMBDA}
.param ln4 = {2*LAMBDA}
.param ln5 = {2*LAMBDA}
.param ln6 = {2*LAMBDA}
.param ln7 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param wp3 = wn1
.param wp4 = wn1
.param wp5 = wn1
.param wp6 = wn1
.param wp7 = wn1 

.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}
.param lp3 = {LAMBDA}
.param lp4 = {LAMBDA}
.param lp5 = {LAMBDA}
.param lp6 = {LAMBDA}
.param lp7 = {LAMBDA}

.global gnd

// inputs 

Vdd vdd gnd 'SUPPLY'


V_in_a0 node_a0 gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_a1 node_a1 gnd PULSE(0 1.8 0ns 100ps 100ps 30ns 50ns)
V_in_a2 node_a2 gnd PULSE(0 1.8 0ns 100ps 100ps 40ns 60ns)
V_in_a3 node_a3 gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)

V_in_b0 node_b0 gnd PULSE(0 1.8 0ns 100ps 100ps 60ns 80ns)
V_in_b1 node_b1 gnd PULSE(0 1.8 0ns 100ps 100ps 70ns 90ns)
V_in_b2 node_b2 gnd PULSE(0 1.8 0ns 100ps 100ps 80ns 100ns)
V_in_b3 node_b3 gnd PULSE(0 1.8 0ns 100ps 100ps 90ns 110ns)

V_in_s0 node_s0 gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 50ns)
V_in_s1 node_s1 gnd PULSE(0 1.8 0ns 100ps 100ps 30ns 60ns)

X1 node_s0 node_s1 node_a0 node_a1 node_a2 node_a3 node_b0 node_b1 node_b2 node_b3 node_sa0 node_sa1 node_sa2 node_sa3 node_sac node_ss0 node_ss1 node_ss2 node_ss3 node_ssc node_cg1 node_ce2 node_cl3 node_r0 node_r1 node_r2 node_r3 vdd gnd alu


C1 node_sa0 gnd 100f
C2 node_sa1 gnd 100f
C3 node_sa2 gnd 100f
C4 node_sa3 gnd 100f
C5 node_sac gnd 100f
C6 node_ss0 gnd 100f
C7 node_ss1 gnd 100f
C8 node_ss2 gnd 100f
C9 node_ss3 gnd 100f
C10 node_ssc gnd 100f
C11 node_cg1 gnd 100f
C12 node_ce2 gnd 100f
C13 node_cl3 gnd 100f
C14 node_r0 gnd 100f
C15 node_r1 gnd 100f
C16 node_r2 gnd 100f
C17 node_r3 gnd 100f


* .tran 1n 1500n

* .control
* run
* set color0 = rgb:f/f/e
* set color1 = black
* plot v(node_s0) v(node_s1)+2 v(node_a0)+4 v(node_a1)+6 v(node_a2)+8 v(node_a3)+10 v(node_b0)+12 v(node_b1)+14 v(node_b2)+16 v(node_b3)+18 v(node_cg1)+20 v(node_ce2)+22 v(node_cl3)+24 
* hardcopy image.ps v(node_s0) v(node_s1)+2 v(node_a0)+4 v(node_a1)+6 v(node_a2)+8 v(node_a3)+10 v(node_b0)+12 v(node_b1)+14 v(node_b2)+16 v(node_b3)+18 v(node_cg1)+20 v(node_ce2)+22 v(node_cl3)+24 
* .end
* .endc


.tran 1n 1500n

.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(node_s0) v(node_s1)+2 v(node_a0)+4 v(node_a1)+6 v(node_a2)+8 v(node_a3)+10 v(node_b0)+12 v(node_b1)+14 v(node_b2)+16 v(node_b3)+18 v(node_sa0)+20 v(node_sa1)+22 v(node_sa2)+24 v(node_sa3)+26 v(node_sac)+28
hardcopy image.ps v(node_s0) v(node_s1)+2 v(node_a0)+4 v(node_a1)+6 v(node_a2)+8 v(node_a3)+10 v(node_b0)+12 v(node_b1)+14 v(node_b2)+16 v(node_b3)+18 v(node_sa0)+20 v(node_sa1)+22 v(node_sa2)+24 v(node_sa3)+26 v(node_sac)+28
.end
.endc

* .tran 1n 1500n

* .control
* run
* set color0 = rgb:f/f/e
* set color1 = black
* plot v(node_s0) v(node_s1)+2 v(node_a0)+4 v(node_a1)+6 v(node_a2)+8 v(node_a3)+10 v(node_b0)+12 v(node_b1)+14 v(node_b2)+16 v(node_b3)+18 v(node_ss0)+20 v(node_ss1)+22 v(node_ss2)+24 v(node_ss3)+26 v(node_ssc)+28
* hardcopy image.ps v(node_s0) v(node_s1)+2 v(node_a0)+4 v(node_a1)+6 v(node_a2)+8 v(node_a3)+10 v(node_b0)+12 v(node_b1)+14 v(node_b2)+16 v(node_b3)+18 v(node_ss0)+20 v(node_ss1)+22 v(node_ss2)+24 v(node_ss3)+26 v(node_ssc)+28
* .end
* .endc

* .tran 1n 800n

* .control
* run
* set color0 = rgb:f/f/e
* set color1 = black
* plot v(node_s0) v(node_s1)+2 v(node_a0)+4 v(node_a1)+6 v(node_a2)+8 v(node_a3)+10 v(node_b0)+12 v(node_b1)+14 v(node_b2)+16 v(node_b3)+18 v(node_r0)+20 v(node_r1)+22 v(node_r2)+24 v(node_r3)+26
* hardcopy image.ps v(node_s0) v(node_s1)+2 v(node_a0)+4 v(node_a1)+6 v(node_a2)+8 v(node_a3)+10 v(node_b0)+12 v(node_b1)+14 v(node_b2)+16 v(node_b3)+18 v(node_r0)+20 v(node_r1)+22 v(node_r2)+24 v(node_r3)+26
* .end
* .endc