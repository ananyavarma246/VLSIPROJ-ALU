magic
tech scmos
timestamp 1699112416
<< nwell >>
rect -594 810 -319 851
<< ntransistor >>
rect -572 726 -568 737
rect -526 726 -522 737
rect -481 726 -477 737
rect -438 726 -434 737
rect -393 726 -389 737
rect -350 726 -346 737
<< ptransistor >>
rect -572 829 -568 840
rect -526 829 -522 840
rect -481 829 -477 840
rect -438 829 -434 840
rect -393 829 -389 840
rect -350 829 -346 840
<< ndiffusion >>
rect -584 733 -572 737
rect -588 726 -572 733
rect -568 733 -552 737
rect -568 726 -548 733
rect -540 733 -526 737
rect -544 726 -526 733
rect -522 733 -508 737
rect -522 726 -504 733
rect -496 733 -481 737
rect -500 726 -481 733
rect -477 733 -464 737
rect -477 726 -460 733
rect -452 733 -438 737
rect -456 726 -438 733
rect -434 733 -420 737
rect -434 726 -416 733
rect -408 733 -393 737
rect -412 726 -393 733
rect -389 733 -376 737
rect -389 726 -372 733
rect -364 733 -350 737
rect -368 726 -350 733
rect -346 733 -332 737
rect -346 726 -328 733
<< pdiffusion >>
rect -584 836 -572 840
rect -588 829 -572 836
rect -568 836 -552 840
rect -568 829 -548 836
rect -540 836 -526 840
rect -544 829 -526 836
rect -522 836 -508 840
rect -522 829 -504 836
rect -496 836 -481 840
rect -500 829 -481 836
rect -477 836 -464 840
rect -477 829 -460 836
rect -452 836 -438 840
rect -456 829 -438 836
rect -434 836 -420 840
rect -434 829 -416 836
rect -408 836 -393 840
rect -412 829 -393 836
rect -389 836 -376 840
rect -389 829 -372 836
rect -364 836 -350 840
rect -368 829 -350 836
rect -346 836 -332 840
rect -346 829 -328 836
<< ndcontact >>
rect -588 733 -584 737
rect -552 733 -548 737
rect -544 733 -540 737
rect -508 733 -504 737
rect -500 733 -496 737
rect -464 733 -460 737
rect -456 733 -452 737
rect -420 733 -416 737
rect -412 733 -408 737
rect -376 733 -372 737
rect -368 733 -364 737
rect -332 733 -328 737
<< pdcontact >>
rect -588 836 -584 840
rect -552 836 -548 840
rect -544 836 -540 840
rect -508 836 -504 840
rect -500 836 -496 840
rect -464 836 -460 840
rect -456 836 -452 840
rect -420 836 -416 840
rect -412 836 -408 840
rect -376 836 -372 840
rect -368 836 -364 840
rect -332 836 -328 840
<< polysilicon >>
rect -572 840 -568 845
rect -526 840 -522 845
rect -481 840 -477 845
rect -438 840 -434 845
rect -393 840 -389 845
rect -350 840 -346 845
rect -572 737 -568 829
rect -526 782 -522 829
rect -527 773 -522 782
rect -481 781 -477 829
rect -438 781 -434 829
rect -526 737 -522 773
rect -479 772 -477 781
rect -436 772 -434 781
rect -393 779 -389 829
rect -481 737 -477 772
rect -438 737 -434 772
rect -392 770 -389 779
rect -393 737 -389 770
rect -350 737 -346 829
rect -572 719 -568 726
rect -526 719 -522 726
rect -481 719 -477 726
rect -438 719 -434 726
rect -393 719 -389 726
rect -350 719 -346 726
<< polycontact >>
rect -581 774 -572 783
rect -536 773 -527 782
rect -488 772 -479 781
rect -445 772 -436 781
rect -401 770 -392 779
rect -360 778 -350 787
<< metal1 >>
rect -595 852 -319 867
rect -588 840 -584 852
rect -544 840 -540 852
rect -500 840 -496 852
rect -456 840 -452 852
rect -412 840 -408 852
rect -368 840 -364 852
rect -552 825 -548 836
rect -508 825 -504 836
rect -464 825 -460 836
rect -420 825 -416 836
rect -376 825 -372 836
rect -552 821 -372 825
rect -376 787 -367 821
rect -332 790 -328 836
rect -590 774 -581 783
rect -545 773 -536 782
rect -497 772 -488 781
rect -454 772 -445 781
rect -410 770 -401 779
rect -376 778 -360 787
rect -332 778 -320 790
rect -376 737 -372 778
rect -332 737 -328 778
rect -548 733 -544 737
rect -504 733 -500 737
rect -460 733 -456 737
rect -416 733 -412 737
rect -588 719 -584 733
rect -368 719 -364 733
rect -591 704 -315 719
<< labels >>
rlabel metal1 -567 858 -567 858 1 vdd
rlabel metal1 -584 777 -584 777 1 node_a
rlabel metal1 -541 777 -541 777 1 node_b
rlabel metal1 -494 776 -494 776 1 node_c
rlabel metal1 -449 776 -449 776 1 node_d
rlabel metal1 -405 774 -405 774 1 node_e
rlabel metal1 -371 784 -371 784 1 node_nand
rlabel metal1 -512 709 -512 709 1 gnd
rlabel metal1 -547 734 -547 734 1 node_x
rlabel metal1 -502 734 -502 734 1 node_y
rlabel metal1 -458 736 -458 736 1 node_n
rlabel metal1 -414 734 -414 734 1 node_m
rlabel metal1 -325 782 -325 782 1 node_out
<< end >>
