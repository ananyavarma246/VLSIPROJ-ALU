.include TSMC_180nm.txt
.include nor.sub

// parameters
.param SUPPLY = 1.8
.param LAMBDA = 0.18u


.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param wn3 = {10*LAMBDA}
.param wn4 = {10*LAMBDA}
.param wn5 = {10*LAMBDA}
.param wn6 = {10*LAMBDA}
.param wn7 = {10*LAMBDA}

.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}
.param ln3 = {2*LAMBDA}
.param ln4 = {2*LAMBDA}
.param ln5 = {2*LAMBDA}
.param ln6 = {2*LAMBDA}
.param ln7 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param wp3 = wn1
.param wp4 = wn1
.param wp5 = wn1
.param wp6 = wn1
.param wp7 = wn1 

.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}
.param lp3 = {LAMBDA}
.param lp4 = {LAMBDA}
.param lp5 = {LAMBDA}
.param lp6 = {LAMBDA}
.param lp7 = {LAMBDA}

.global gnd


Vdd node_x gnd 'SUPPLY'

V_in_a node_a gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 50ns)
V_in_b node_b gnd PULSE(0 1.8 0ns 100ps 100ps 30ns 60ns)

X1 node_a node_b node_out node_x gnd nor

C1 node_out gnd 100f


.tran 1n 800n

.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(node_a) v(node_b)+2 v(node_out)+4
hardcopy image.ps v(node_a) v(node_b)+2 v(node_out)+4
.end
.endc