magic
tech scmos
timestamp 1701457681
<< nwell >>
rect 488 2020 676 2059
rect 706 2020 894 2059
rect 939 2022 1127 2061
rect 1199 2023 1387 2062
rect 517 1822 705 1861
rect 744 1822 844 1852
rect 917 1808 987 1824
rect 1143 1819 1331 1858
rect 1370 1819 1470 1849
rect 1543 1805 1613 1821
rect 1743 1819 1931 1858
rect 1970 1819 2070 1849
rect 2346 1822 2534 1861
rect 2573 1822 2673 1852
rect 2143 1805 2213 1821
rect 2746 1808 2816 1824
rect 760 1683 860 1713
rect 1386 1680 1486 1710
rect 1986 1680 2086 1710
rect 2589 1683 2689 1713
rect 527 1566 715 1605
rect 1153 1563 1341 1602
rect 1753 1563 1941 1602
rect 2356 1566 2544 1605
rect 541 1205 729 1244
rect 759 1205 947 1244
rect 992 1207 1180 1246
rect 1252 1208 1440 1247
rect -88 1087 -75 1092
rect -359 1085 -346 1086
rect -416 1055 -316 1085
rect -280 1056 -180 1086
rect -145 1057 -45 1087
rect 49 1085 62 1090
rect -8 1055 92 1085
rect 570 1007 758 1046
rect 797 1007 897 1037
rect 970 993 1040 1009
rect 1196 1004 1384 1043
rect 1423 1004 1523 1034
rect 1596 990 1666 1006
rect 1796 1004 1984 1043
rect 2023 1004 2123 1034
rect 2399 1007 2587 1046
rect 2626 1007 2726 1037
rect 2196 990 2266 1006
rect 2799 993 2869 1009
rect -360 965 -347 970
rect -214 966 -201 971
rect -84 969 -71 974
rect -417 935 -317 965
rect -271 936 -171 966
rect -141 939 -41 969
rect 57 968 70 973
rect 0 938 100 968
rect 813 868 913 898
rect 1439 865 1539 895
rect 2039 865 2139 895
rect 2642 868 2742 898
rect 580 751 768 790
rect 1206 748 1394 787
rect 1806 748 1994 787
rect 2409 751 2597 790
rect -69 644 -56 649
rect -340 642 -327 643
rect -397 612 -297 642
rect -261 613 -161 643
rect -126 614 -26 644
rect 68 642 81 647
rect 11 612 111 642
rect -341 522 -328 527
rect -195 523 -182 528
rect -65 526 -52 531
rect -398 492 -298 522
rect -252 493 -152 523
rect -122 496 -22 526
rect 76 525 89 530
rect 19 495 119 525
rect -1058 438 -958 468
rect -1249 414 -1174 436
rect -1056 337 -956 367
rect -1053 238 -953 268
rect -56 219 -43 224
rect -327 217 -314 218
rect -1251 195 -1176 217
rect -384 187 -284 217
rect -248 188 -148 218
rect -113 189 -13 219
rect 81 217 94 222
rect 24 187 124 217
rect -1051 130 -951 160
rect -328 97 -315 102
rect -182 98 -169 103
rect -52 101 -39 106
rect -385 67 -285 97
rect -239 68 -139 98
rect -109 71 -9 101
rect 89 100 102 105
rect 32 70 132 100
rect 2067 -2 2142 20
rect 2337 -7 2412 15
rect 2592 -1 2667 21
rect 2860 -1 2935 21
rect 3419 -156 3597 -121
rect 2213 -213 2488 -172
rect 2595 -213 2870 -172
rect 2977 -213 3252 -172
rect -4 -231 9 -226
rect -275 -233 -262 -232
rect -332 -263 -232 -233
rect -196 -262 -96 -232
rect -61 -261 39 -231
rect 133 -233 146 -228
rect 76 -263 176 -233
rect 2035 -275 2135 -245
rect -276 -353 -263 -348
rect -130 -352 -117 -347
rect 0 -349 13 -344
rect -333 -383 -233 -353
rect -187 -382 -87 -352
rect -57 -379 43 -349
rect 141 -350 154 -345
rect 84 -380 184 -350
rect 395 -443 495 -413
rect -276 -549 -176 -519
rect 2051 -530 2255 -498
rect -100 -605 0 -575
rect 154 -615 254 -585
rect 2050 -777 2254 -745
rect 2404 -833 2679 -792
rect 2054 -1003 2258 -971
rect 2051 -1210 2255 -1178
rect 2078 -1420 2178 -1390
rect 2264 -1439 2539 -1398
rect 2636 -1438 2911 -1397
rect 3010 -1438 3285 -1397
rect 3469 -1483 3647 -1448
rect 2094 -1541 2169 -1519
rect 2291 -1587 2366 -1565
rect 2699 -1611 2774 -1589
rect 3126 -1610 3201 -1588
<< ntransistor >>
rect 503 1962 506 1969
rect 532 1962 534 1969
rect 563 1962 566 1969
rect 592 1962 595 1969
rect 621 1962 624 1969
rect 651 1962 654 1969
rect 721 1962 724 1969
rect 750 1962 752 1969
rect 781 1962 784 1969
rect 810 1962 813 1969
rect 839 1962 842 1969
rect 869 1962 872 1969
rect 954 1964 957 1971
rect 983 1964 985 1971
rect 1014 1964 1017 1971
rect 1043 1964 1046 1971
rect 1072 1964 1075 1971
rect 1102 1964 1105 1971
rect 1214 1965 1217 1972
rect 1243 1965 1245 1972
rect 1274 1965 1277 1972
rect 1303 1965 1306 1972
rect 1332 1965 1335 1972
rect 1362 1965 1365 1972
rect 759 1776 763 1785
rect 791 1776 795 1785
rect 825 1776 829 1785
rect 932 1773 934 1777
rect 950 1773 952 1777
rect 969 1773 971 1777
rect 532 1764 535 1771
rect 561 1764 563 1771
rect 592 1764 595 1771
rect 621 1764 624 1771
rect 650 1764 653 1771
rect 680 1764 683 1771
rect 1385 1773 1389 1782
rect 1417 1773 1421 1782
rect 1451 1773 1455 1782
rect 1558 1770 1560 1774
rect 1576 1770 1578 1774
rect 1595 1770 1597 1774
rect 1158 1761 1161 1768
rect 1187 1761 1189 1768
rect 1218 1761 1221 1768
rect 1247 1761 1250 1768
rect 1276 1761 1279 1768
rect 1306 1761 1309 1768
rect 1985 1773 1989 1782
rect 2017 1773 2021 1782
rect 2051 1773 2055 1782
rect 2158 1770 2160 1774
rect 2176 1770 2178 1774
rect 2195 1770 2197 1774
rect 2588 1776 2592 1785
rect 2620 1776 2624 1785
rect 2654 1776 2658 1785
rect 2761 1773 2763 1777
rect 2779 1773 2781 1777
rect 2798 1773 2800 1777
rect 1758 1761 1761 1768
rect 1787 1761 1789 1768
rect 1818 1761 1821 1768
rect 1847 1761 1850 1768
rect 1876 1761 1879 1768
rect 1906 1761 1909 1768
rect 2361 1764 2364 1771
rect 2390 1764 2392 1771
rect 2421 1764 2424 1771
rect 2450 1764 2453 1771
rect 2479 1764 2482 1771
rect 2509 1764 2512 1771
rect 775 1637 779 1646
rect 807 1637 811 1646
rect 841 1637 845 1646
rect 1401 1634 1405 1643
rect 1433 1634 1437 1643
rect 1467 1634 1471 1643
rect 2001 1634 2005 1643
rect 2033 1634 2037 1643
rect 2067 1634 2071 1643
rect 2604 1637 2608 1646
rect 2636 1637 2640 1646
rect 2670 1637 2674 1646
rect 542 1508 545 1515
rect 571 1508 573 1515
rect 602 1508 605 1515
rect 631 1508 634 1515
rect 660 1508 663 1515
rect 690 1508 693 1515
rect 1168 1505 1171 1512
rect 1197 1505 1199 1512
rect 1228 1505 1231 1512
rect 1257 1505 1260 1512
rect 1286 1505 1289 1512
rect 1316 1505 1319 1512
rect 1768 1505 1771 1512
rect 1797 1505 1799 1512
rect 1828 1505 1831 1512
rect 1857 1505 1860 1512
rect 1886 1505 1889 1512
rect 1916 1505 1919 1512
rect 2371 1508 2374 1515
rect 2400 1508 2402 1515
rect 2431 1508 2434 1515
rect 2460 1508 2463 1515
rect 2489 1508 2492 1515
rect 2519 1508 2522 1515
rect 556 1147 559 1154
rect 585 1147 587 1154
rect 616 1147 619 1154
rect 645 1147 648 1154
rect 674 1147 677 1154
rect 704 1147 707 1154
rect 774 1147 777 1154
rect 803 1147 805 1154
rect 834 1147 837 1154
rect 863 1147 866 1154
rect 892 1147 895 1154
rect 922 1147 925 1154
rect 1007 1149 1010 1156
rect 1036 1149 1038 1156
rect 1067 1149 1070 1156
rect 1096 1149 1099 1156
rect 1125 1149 1128 1156
rect 1155 1149 1158 1156
rect 1267 1150 1270 1157
rect 1296 1150 1298 1157
rect 1327 1150 1330 1157
rect 1356 1150 1359 1157
rect 1385 1150 1388 1157
rect 1415 1150 1418 1157
rect -401 1009 -397 1018
rect -369 1009 -365 1018
rect -335 1009 -331 1018
rect -265 1010 -261 1019
rect -233 1010 -229 1019
rect -199 1010 -195 1019
rect -130 1011 -126 1020
rect -98 1011 -94 1020
rect -64 1011 -60 1020
rect 7 1009 11 1018
rect 39 1009 43 1018
rect 73 1009 77 1018
rect 812 961 816 970
rect 844 961 848 970
rect 878 961 882 970
rect 985 958 987 962
rect 1003 958 1005 962
rect 1022 958 1024 962
rect -402 889 -398 898
rect -370 889 -366 898
rect -336 889 -332 898
rect -256 890 -252 899
rect -224 890 -220 899
rect -190 890 -186 899
rect -126 893 -122 902
rect -94 893 -90 902
rect -60 893 -56 902
rect 585 949 588 956
rect 614 949 616 956
rect 645 949 648 956
rect 674 949 677 956
rect 703 949 706 956
rect 733 949 736 956
rect 1438 958 1442 967
rect 1470 958 1474 967
rect 1504 958 1508 967
rect 1611 955 1613 959
rect 1629 955 1631 959
rect 1648 955 1650 959
rect 1211 946 1214 953
rect 1240 946 1242 953
rect 1271 946 1274 953
rect 1300 946 1303 953
rect 1329 946 1332 953
rect 1359 946 1362 953
rect 2038 958 2042 967
rect 2070 958 2074 967
rect 2104 958 2108 967
rect 2211 955 2213 959
rect 2229 955 2231 959
rect 2248 955 2250 959
rect 2641 961 2645 970
rect 2673 961 2677 970
rect 2707 961 2711 970
rect 2814 958 2816 962
rect 2832 958 2834 962
rect 2851 958 2853 962
rect 1811 946 1814 953
rect 1840 946 1842 953
rect 1871 946 1874 953
rect 1900 946 1903 953
rect 1929 946 1932 953
rect 1959 946 1962 953
rect 2414 949 2417 956
rect 2443 949 2445 956
rect 2474 949 2477 956
rect 2503 949 2506 956
rect 2532 949 2535 956
rect 2562 949 2565 956
rect 15 892 19 901
rect 47 892 51 901
rect 81 892 85 901
rect 828 822 832 831
rect 860 822 864 831
rect 894 822 898 831
rect 1454 819 1458 828
rect 1486 819 1490 828
rect 1520 819 1524 828
rect 2054 819 2058 828
rect 2086 819 2090 828
rect 2120 819 2124 828
rect 2657 822 2661 831
rect 2689 822 2693 831
rect 2723 822 2727 831
rect 595 693 598 700
rect 624 693 626 700
rect 655 693 658 700
rect 684 693 687 700
rect 713 693 716 700
rect 743 693 746 700
rect 1221 690 1224 697
rect 1250 690 1252 697
rect 1281 690 1284 697
rect 1310 690 1313 697
rect 1339 690 1342 697
rect 1369 690 1372 697
rect 1821 690 1824 697
rect 1850 690 1852 697
rect 1881 690 1884 697
rect 1910 690 1913 697
rect 1939 690 1942 697
rect 1969 690 1972 697
rect 2424 693 2427 700
rect 2453 693 2455 700
rect 2484 693 2487 700
rect 2513 693 2516 700
rect 2542 693 2545 700
rect 2572 693 2575 700
rect -382 566 -378 575
rect -350 566 -346 575
rect -316 566 -312 575
rect -246 567 -242 576
rect -214 567 -210 576
rect -180 567 -176 576
rect -111 568 -107 577
rect -79 568 -75 577
rect -45 568 -41 577
rect 26 566 30 575
rect 58 566 62 575
rect 92 566 96 575
rect -383 446 -379 455
rect -351 446 -347 455
rect -317 446 -313 455
rect -237 447 -233 456
rect -205 447 -201 456
rect -171 447 -167 456
rect -107 450 -103 459
rect -75 450 -71 459
rect -41 450 -37 459
rect 34 449 38 458
rect 66 449 70 458
rect 100 449 104 458
rect -1043 392 -1039 401
rect -1011 392 -1007 401
rect -977 392 -973 401
rect -1215 378 -1211 392
rect -1041 291 -1037 300
rect -1009 291 -1005 300
rect -975 291 -971 300
rect -1038 192 -1034 201
rect -1006 192 -1002 201
rect -972 192 -968 201
rect -1217 159 -1213 173
rect -369 141 -365 150
rect -337 141 -333 150
rect -303 141 -299 150
rect -233 142 -229 151
rect -201 142 -197 151
rect -167 142 -163 151
rect -98 143 -94 152
rect -66 143 -62 152
rect -32 143 -28 152
rect 39 141 43 150
rect 71 141 75 150
rect 105 141 109 150
rect -1036 84 -1032 93
rect -1004 84 -1000 93
rect -970 84 -966 93
rect -370 21 -366 30
rect -338 21 -334 30
rect -304 21 -300 30
rect -224 22 -220 31
rect -192 22 -188 31
rect -158 22 -154 31
rect -94 25 -90 34
rect -62 25 -58 34
rect -28 25 -24 34
rect 47 24 51 33
rect 79 24 83 33
rect 113 24 117 33
rect 2101 -38 2105 -24
rect 2371 -43 2375 -29
rect 2626 -37 2630 -23
rect 2894 -37 2898 -23
rect -317 -309 -313 -300
rect -285 -309 -281 -300
rect -251 -309 -247 -300
rect -181 -308 -177 -299
rect -149 -308 -145 -299
rect -115 -308 -111 -299
rect -46 -307 -42 -298
rect -14 -307 -10 -298
rect 20 -307 24 -298
rect 91 -309 95 -300
rect 123 -309 127 -300
rect 157 -309 161 -300
rect 3438 -224 3442 -215
rect 3473 -224 3477 -215
rect 3506 -224 3510 -215
rect 3539 -224 3543 -215
rect 3572 -224 3576 -215
rect 2235 -297 2239 -286
rect 2281 -297 2285 -286
rect 2326 -297 2330 -286
rect 2369 -297 2373 -286
rect 2414 -297 2418 -286
rect 2457 -297 2461 -286
rect 2617 -297 2621 -286
rect 2663 -297 2667 -286
rect 2708 -297 2712 -286
rect 2751 -297 2755 -286
rect 2796 -297 2800 -286
rect 2839 -297 2843 -286
rect 2999 -297 3003 -286
rect 3045 -297 3049 -286
rect 3090 -297 3094 -286
rect 3133 -297 3137 -286
rect 3178 -297 3182 -286
rect 3221 -297 3225 -286
rect 2050 -321 2054 -312
rect 2082 -321 2086 -312
rect 2116 -321 2120 -312
rect -318 -429 -314 -420
rect -286 -429 -282 -420
rect -252 -429 -248 -420
rect -172 -428 -168 -419
rect -140 -428 -136 -419
rect -106 -428 -102 -419
rect -42 -425 -38 -416
rect -10 -425 -6 -416
rect 24 -425 28 -416
rect 99 -426 103 -417
rect 131 -426 135 -417
rect 165 -426 169 -417
rect 410 -489 414 -480
rect 442 -489 446 -480
rect 476 -489 480 -480
rect -261 -595 -257 -586
rect -229 -595 -225 -586
rect -195 -595 -191 -586
rect -85 -651 -81 -642
rect -53 -651 -49 -642
rect -19 -651 -15 -642
rect 2067 -605 2070 -599
rect 2102 -605 2105 -599
rect 2137 -605 2140 -599
rect 2169 -605 2172 -599
rect 2200 -605 2203 -599
rect 2233 -605 2236 -599
rect 169 -661 173 -652
rect 201 -661 205 -652
rect 235 -661 239 -652
rect 2066 -852 2069 -846
rect 2101 -852 2104 -846
rect 2136 -852 2139 -846
rect 2168 -852 2171 -846
rect 2199 -852 2202 -846
rect 2232 -852 2235 -846
rect 2426 -917 2430 -906
rect 2472 -917 2476 -906
rect 2517 -917 2521 -906
rect 2560 -917 2564 -906
rect 2605 -917 2609 -906
rect 2648 -917 2652 -906
rect 2070 -1078 2073 -1072
rect 2105 -1078 2108 -1072
rect 2140 -1078 2143 -1072
rect 2172 -1078 2175 -1072
rect 2203 -1078 2206 -1072
rect 2236 -1078 2239 -1072
rect 2067 -1285 2070 -1279
rect 2102 -1285 2105 -1279
rect 2137 -1285 2140 -1279
rect 2169 -1285 2172 -1279
rect 2200 -1285 2203 -1279
rect 2233 -1285 2236 -1279
rect 2093 -1466 2097 -1457
rect 2125 -1466 2129 -1457
rect 2159 -1466 2163 -1457
rect 2286 -1523 2290 -1512
rect 2332 -1523 2336 -1512
rect 2377 -1523 2381 -1512
rect 2420 -1523 2424 -1512
rect 2465 -1523 2469 -1512
rect 2508 -1523 2512 -1512
rect 2658 -1522 2662 -1511
rect 2704 -1522 2708 -1511
rect 2749 -1522 2753 -1511
rect 2792 -1522 2796 -1511
rect 2837 -1522 2841 -1511
rect 2880 -1522 2884 -1511
rect 3032 -1522 3036 -1511
rect 3078 -1522 3082 -1511
rect 3123 -1522 3127 -1511
rect 3166 -1522 3170 -1511
rect 3211 -1522 3215 -1511
rect 3254 -1522 3258 -1511
rect 3488 -1551 3492 -1542
rect 3523 -1551 3527 -1542
rect 3556 -1551 3560 -1542
rect 3589 -1551 3593 -1542
rect 3622 -1551 3626 -1542
rect 2128 -1577 2132 -1563
rect 2325 -1623 2329 -1609
rect 2733 -1647 2737 -1633
rect 3160 -1646 3164 -1632
<< ptransistor >>
rect 503 2034 506 2041
rect 532 2034 534 2041
rect 563 2034 566 2041
rect 592 2034 595 2041
rect 621 2034 624 2041
rect 651 2034 654 2041
rect 721 2034 724 2041
rect 750 2034 752 2041
rect 781 2034 784 2041
rect 810 2034 813 2041
rect 839 2034 842 2041
rect 869 2034 872 2041
rect 954 2036 957 2043
rect 983 2036 985 2043
rect 1014 2036 1017 2043
rect 1043 2036 1046 2043
rect 1072 2036 1075 2043
rect 1102 2036 1105 2043
rect 1214 2037 1217 2044
rect 1243 2037 1245 2044
rect 1274 2037 1277 2044
rect 1303 2037 1306 2044
rect 1332 2037 1335 2044
rect 1362 2037 1365 2044
rect 532 1836 535 1843
rect 561 1836 563 1843
rect 592 1836 595 1843
rect 621 1836 624 1843
rect 650 1836 653 1843
rect 680 1836 683 1843
rect 759 1834 763 1843
rect 791 1834 795 1843
rect 825 1834 829 1843
rect 1158 1833 1161 1840
rect 1187 1833 1189 1840
rect 1218 1833 1221 1840
rect 1247 1833 1250 1840
rect 1276 1833 1279 1840
rect 1306 1833 1309 1840
rect 932 1814 934 1818
rect 950 1814 952 1818
rect 969 1814 971 1818
rect 1385 1831 1389 1840
rect 1417 1831 1421 1840
rect 1451 1831 1455 1840
rect 1758 1833 1761 1840
rect 1787 1833 1789 1840
rect 1818 1833 1821 1840
rect 1847 1833 1850 1840
rect 1876 1833 1879 1840
rect 1906 1833 1909 1840
rect 1558 1811 1560 1815
rect 1576 1811 1578 1815
rect 1595 1811 1597 1815
rect 1985 1831 1989 1840
rect 2017 1831 2021 1840
rect 2051 1831 2055 1840
rect 2361 1836 2364 1843
rect 2390 1836 2392 1843
rect 2421 1836 2424 1843
rect 2450 1836 2453 1843
rect 2479 1836 2482 1843
rect 2509 1836 2512 1843
rect 2158 1811 2160 1815
rect 2176 1811 2178 1815
rect 2195 1811 2197 1815
rect 2588 1834 2592 1843
rect 2620 1834 2624 1843
rect 2654 1834 2658 1843
rect 2761 1814 2763 1818
rect 2779 1814 2781 1818
rect 2798 1814 2800 1818
rect 775 1695 779 1704
rect 807 1695 811 1704
rect 841 1695 845 1704
rect 1401 1692 1405 1701
rect 1433 1692 1437 1701
rect 1467 1692 1471 1701
rect 2001 1692 2005 1701
rect 2033 1692 2037 1701
rect 2067 1692 2071 1701
rect 2604 1695 2608 1704
rect 2636 1695 2640 1704
rect 2670 1695 2674 1704
rect 542 1580 545 1587
rect 571 1580 573 1587
rect 602 1580 605 1587
rect 631 1580 634 1587
rect 660 1580 663 1587
rect 690 1580 693 1587
rect 1168 1577 1171 1584
rect 1197 1577 1199 1584
rect 1228 1577 1231 1584
rect 1257 1577 1260 1584
rect 1286 1577 1289 1584
rect 1316 1577 1319 1584
rect 1768 1577 1771 1584
rect 1797 1577 1799 1584
rect 1828 1577 1831 1584
rect 1857 1577 1860 1584
rect 1886 1577 1889 1584
rect 1916 1577 1919 1584
rect 2371 1580 2374 1587
rect 2400 1580 2402 1587
rect 2431 1580 2434 1587
rect 2460 1580 2463 1587
rect 2489 1580 2492 1587
rect 2519 1580 2522 1587
rect 556 1219 559 1226
rect 585 1219 587 1226
rect 616 1219 619 1226
rect 645 1219 648 1226
rect 674 1219 677 1226
rect 704 1219 707 1226
rect 774 1219 777 1226
rect 803 1219 805 1226
rect 834 1219 837 1226
rect 863 1219 866 1226
rect 892 1219 895 1226
rect 922 1219 925 1226
rect 1007 1221 1010 1228
rect 1036 1221 1038 1228
rect 1067 1221 1070 1228
rect 1096 1221 1099 1228
rect 1125 1221 1128 1228
rect 1155 1221 1158 1228
rect 1267 1222 1270 1229
rect 1296 1222 1298 1229
rect 1327 1222 1330 1229
rect 1356 1222 1359 1229
rect 1385 1222 1388 1229
rect 1415 1222 1418 1229
rect -401 1067 -397 1076
rect -369 1067 -365 1076
rect -335 1067 -331 1076
rect -265 1068 -261 1077
rect -233 1068 -229 1077
rect -199 1068 -195 1077
rect -130 1069 -126 1078
rect -98 1069 -94 1078
rect -64 1069 -60 1078
rect 7 1067 11 1076
rect 39 1067 43 1076
rect 73 1067 77 1076
rect 585 1021 588 1028
rect 614 1021 616 1028
rect 645 1021 648 1028
rect 674 1021 677 1028
rect 703 1021 706 1028
rect 733 1021 736 1028
rect -402 947 -398 956
rect -370 947 -366 956
rect -336 947 -332 956
rect -256 948 -252 957
rect -224 948 -220 957
rect -190 948 -186 957
rect -126 951 -122 960
rect -94 951 -90 960
rect -60 951 -56 960
rect 15 950 19 959
rect 47 950 51 959
rect 81 950 85 959
rect 812 1019 816 1028
rect 844 1019 848 1028
rect 878 1019 882 1028
rect 1211 1018 1214 1025
rect 1240 1018 1242 1025
rect 1271 1018 1274 1025
rect 1300 1018 1303 1025
rect 1329 1018 1332 1025
rect 1359 1018 1362 1025
rect 985 999 987 1003
rect 1003 999 1005 1003
rect 1022 999 1024 1003
rect 1438 1016 1442 1025
rect 1470 1016 1474 1025
rect 1504 1016 1508 1025
rect 1811 1018 1814 1025
rect 1840 1018 1842 1025
rect 1871 1018 1874 1025
rect 1900 1018 1903 1025
rect 1929 1018 1932 1025
rect 1959 1018 1962 1025
rect 1611 996 1613 1000
rect 1629 996 1631 1000
rect 1648 996 1650 1000
rect 2038 1016 2042 1025
rect 2070 1016 2074 1025
rect 2104 1016 2108 1025
rect 2414 1021 2417 1028
rect 2443 1021 2445 1028
rect 2474 1021 2477 1028
rect 2503 1021 2506 1028
rect 2532 1021 2535 1028
rect 2562 1021 2565 1028
rect 2211 996 2213 1000
rect 2229 996 2231 1000
rect 2248 996 2250 1000
rect 2641 1019 2645 1028
rect 2673 1019 2677 1028
rect 2707 1019 2711 1028
rect 2814 999 2816 1003
rect 2832 999 2834 1003
rect 2851 999 2853 1003
rect 828 880 832 889
rect 860 880 864 889
rect 894 880 898 889
rect 1454 877 1458 886
rect 1486 877 1490 886
rect 1520 877 1524 886
rect 2054 877 2058 886
rect 2086 877 2090 886
rect 2120 877 2124 886
rect 2657 880 2661 889
rect 2689 880 2693 889
rect 2723 880 2727 889
rect 595 765 598 772
rect 624 765 626 772
rect 655 765 658 772
rect 684 765 687 772
rect 713 765 716 772
rect 743 765 746 772
rect 1221 762 1224 769
rect 1250 762 1252 769
rect 1281 762 1284 769
rect 1310 762 1313 769
rect 1339 762 1342 769
rect 1369 762 1372 769
rect 1821 762 1824 769
rect 1850 762 1852 769
rect 1881 762 1884 769
rect 1910 762 1913 769
rect 1939 762 1942 769
rect 1969 762 1972 769
rect 2424 765 2427 772
rect 2453 765 2455 772
rect 2484 765 2487 772
rect 2513 765 2516 772
rect 2542 765 2545 772
rect 2572 765 2575 772
rect -382 624 -378 633
rect -350 624 -346 633
rect -316 624 -312 633
rect -246 625 -242 634
rect -214 625 -210 634
rect -180 625 -176 634
rect -111 626 -107 635
rect -79 626 -75 635
rect -45 626 -41 635
rect 26 624 30 633
rect 58 624 62 633
rect 92 624 96 633
rect -383 504 -379 513
rect -351 504 -347 513
rect -317 504 -313 513
rect -237 505 -233 514
rect -205 505 -201 514
rect -171 505 -167 514
rect -107 508 -103 517
rect -75 508 -71 517
rect -41 508 -37 517
rect -1043 450 -1039 459
rect -1011 450 -1007 459
rect -977 450 -973 459
rect 34 507 38 516
rect 66 507 70 516
rect 100 507 104 516
rect -1215 420 -1211 430
rect -1041 349 -1037 358
rect -1009 349 -1005 358
rect -975 349 -971 358
rect -1038 250 -1034 259
rect -1006 250 -1002 259
rect -972 250 -968 259
rect -1217 201 -1213 211
rect -369 199 -365 208
rect -337 199 -333 208
rect -303 199 -299 208
rect -233 200 -229 209
rect -201 200 -197 209
rect -167 200 -163 209
rect -98 201 -94 210
rect -66 201 -62 210
rect -32 201 -28 210
rect -1036 142 -1032 151
rect -1004 142 -1000 151
rect -970 142 -966 151
rect 39 199 43 208
rect 71 199 75 208
rect 105 199 109 208
rect -370 79 -366 88
rect -338 79 -334 88
rect -304 79 -300 88
rect -224 80 -220 89
rect -192 80 -188 89
rect -158 80 -154 89
rect -94 83 -90 92
rect -62 83 -58 92
rect -28 83 -24 92
rect 47 82 51 91
rect 79 82 83 91
rect 113 82 117 91
rect 2101 4 2105 14
rect 2371 -1 2375 9
rect 2626 5 2630 15
rect 2894 5 2898 15
rect 3438 -142 3442 -133
rect 3473 -142 3477 -133
rect 3506 -142 3510 -133
rect 3539 -142 3543 -133
rect 3572 -142 3576 -133
rect 2235 -194 2239 -183
rect 2281 -194 2285 -183
rect 2326 -194 2330 -183
rect 2369 -194 2373 -183
rect 2414 -194 2418 -183
rect 2457 -194 2461 -183
rect 2617 -194 2621 -183
rect 2663 -194 2667 -183
rect 2708 -194 2712 -183
rect 2751 -194 2755 -183
rect 2796 -194 2800 -183
rect 2839 -194 2843 -183
rect 2999 -194 3003 -183
rect 3045 -194 3049 -183
rect 3090 -194 3094 -183
rect 3133 -194 3137 -183
rect 3178 -194 3182 -183
rect 3221 -194 3225 -183
rect -317 -251 -313 -242
rect -285 -251 -281 -242
rect -251 -251 -247 -242
rect -181 -250 -177 -241
rect -149 -250 -145 -241
rect -115 -250 -111 -241
rect -46 -249 -42 -240
rect -14 -249 -10 -240
rect 20 -249 24 -240
rect 91 -251 95 -242
rect 123 -251 127 -242
rect 157 -251 161 -242
rect 2050 -263 2054 -254
rect 2082 -263 2086 -254
rect 2116 -263 2120 -254
rect -318 -371 -314 -362
rect -286 -371 -282 -362
rect -252 -371 -248 -362
rect -172 -370 -168 -361
rect -140 -370 -136 -361
rect -106 -370 -102 -361
rect -42 -367 -38 -358
rect -10 -367 -6 -358
rect 24 -367 28 -358
rect 99 -368 103 -359
rect 131 -368 135 -359
rect 165 -368 169 -359
rect 410 -431 414 -422
rect 442 -431 446 -422
rect 476 -431 480 -422
rect 2067 -516 2070 -510
rect 2102 -516 2105 -510
rect 2137 -516 2140 -510
rect 2169 -516 2172 -510
rect 2200 -516 2203 -510
rect 2233 -516 2236 -510
rect -261 -537 -257 -528
rect -229 -537 -225 -528
rect -195 -537 -191 -528
rect -85 -593 -81 -584
rect -53 -593 -49 -584
rect -19 -593 -15 -584
rect 169 -603 173 -594
rect 201 -603 205 -594
rect 235 -603 239 -594
rect 2066 -763 2069 -757
rect 2101 -763 2104 -757
rect 2136 -763 2139 -757
rect 2168 -763 2171 -757
rect 2199 -763 2202 -757
rect 2232 -763 2235 -757
rect 2426 -814 2430 -803
rect 2472 -814 2476 -803
rect 2517 -814 2521 -803
rect 2560 -814 2564 -803
rect 2605 -814 2609 -803
rect 2648 -814 2652 -803
rect 2070 -989 2073 -983
rect 2105 -989 2108 -983
rect 2140 -989 2143 -983
rect 2172 -989 2175 -983
rect 2203 -989 2206 -983
rect 2236 -989 2239 -983
rect 2067 -1196 2070 -1190
rect 2102 -1196 2105 -1190
rect 2137 -1196 2140 -1190
rect 2169 -1196 2172 -1190
rect 2200 -1196 2203 -1190
rect 2233 -1196 2236 -1190
rect 2093 -1408 2097 -1399
rect 2125 -1408 2129 -1399
rect 2159 -1408 2163 -1399
rect 2286 -1420 2290 -1409
rect 2332 -1420 2336 -1409
rect 2377 -1420 2381 -1409
rect 2420 -1420 2424 -1409
rect 2465 -1420 2469 -1409
rect 2508 -1420 2512 -1409
rect 2658 -1419 2662 -1408
rect 2704 -1419 2708 -1408
rect 2749 -1419 2753 -1408
rect 2792 -1419 2796 -1408
rect 2837 -1419 2841 -1408
rect 2880 -1419 2884 -1408
rect 3032 -1419 3036 -1408
rect 3078 -1419 3082 -1408
rect 3123 -1419 3127 -1408
rect 3166 -1419 3170 -1408
rect 3211 -1419 3215 -1408
rect 3254 -1419 3258 -1408
rect 3488 -1469 3492 -1460
rect 3523 -1469 3527 -1460
rect 3556 -1469 3560 -1460
rect 3589 -1469 3593 -1460
rect 3622 -1469 3626 -1460
rect 2128 -1535 2132 -1525
rect 2325 -1581 2329 -1571
rect 2733 -1605 2737 -1595
rect 3160 -1604 3164 -1594
<< ndiffusion >>
rect 498 1965 503 1969
rect 494 1962 503 1965
rect 506 1965 515 1969
rect 506 1962 519 1965
rect 527 1965 532 1969
rect 523 1962 532 1965
rect 534 1965 544 1969
rect 534 1962 548 1965
rect 556 1965 563 1969
rect 552 1962 563 1965
rect 566 1965 573 1969
rect 566 1962 577 1965
rect 585 1965 592 1969
rect 581 1962 592 1965
rect 595 1965 602 1969
rect 595 1962 606 1965
rect 614 1965 621 1969
rect 610 1962 621 1965
rect 624 1965 631 1969
rect 624 1962 635 1965
rect 643 1965 651 1969
rect 639 1962 651 1965
rect 654 1965 660 1969
rect 654 1962 664 1965
rect 716 1965 721 1969
rect 712 1962 721 1965
rect 724 1965 733 1969
rect 724 1962 737 1965
rect 745 1965 750 1969
rect 741 1962 750 1965
rect 752 1965 762 1969
rect 752 1962 766 1965
rect 774 1965 781 1969
rect 770 1962 781 1965
rect 784 1965 791 1969
rect 784 1962 795 1965
rect 803 1965 810 1969
rect 799 1962 810 1965
rect 813 1965 820 1969
rect 813 1962 824 1965
rect 832 1965 839 1969
rect 828 1962 839 1965
rect 842 1965 849 1969
rect 842 1962 853 1965
rect 861 1965 869 1969
rect 857 1962 869 1965
rect 872 1965 878 1969
rect 872 1962 882 1965
rect 949 1967 954 1971
rect 945 1964 954 1967
rect 957 1967 966 1971
rect 957 1964 970 1967
rect 978 1967 983 1971
rect 974 1964 983 1967
rect 985 1967 995 1971
rect 985 1964 999 1967
rect 1007 1967 1014 1971
rect 1003 1964 1014 1967
rect 1017 1967 1024 1971
rect 1017 1964 1028 1967
rect 1036 1967 1043 1971
rect 1032 1964 1043 1967
rect 1046 1967 1053 1971
rect 1046 1964 1057 1967
rect 1065 1967 1072 1971
rect 1061 1964 1072 1967
rect 1075 1967 1082 1971
rect 1075 1964 1086 1967
rect 1094 1967 1102 1971
rect 1090 1964 1102 1967
rect 1105 1967 1111 1971
rect 1105 1964 1115 1967
rect 1209 1968 1214 1972
rect 1205 1965 1214 1968
rect 1217 1968 1226 1972
rect 1217 1965 1230 1968
rect 1238 1968 1243 1972
rect 1234 1965 1243 1968
rect 1245 1968 1255 1972
rect 1245 1965 1259 1968
rect 1267 1968 1274 1972
rect 1263 1965 1274 1968
rect 1277 1968 1284 1972
rect 1277 1965 1288 1968
rect 1296 1968 1303 1972
rect 1292 1965 1303 1968
rect 1306 1968 1313 1972
rect 1306 1965 1317 1968
rect 1325 1968 1332 1972
rect 1321 1965 1332 1968
rect 1335 1968 1342 1972
rect 1335 1965 1346 1968
rect 1354 1968 1362 1972
rect 1350 1965 1362 1968
rect 1365 1968 1371 1972
rect 1365 1965 1375 1968
rect 755 1780 759 1785
rect 750 1776 759 1780
rect 763 1780 769 1785
rect 763 1776 774 1780
rect 786 1780 791 1785
rect 781 1776 791 1780
rect 795 1780 800 1785
rect 795 1776 805 1780
rect 819 1780 825 1785
rect 814 1776 825 1780
rect 829 1780 833 1785
rect 829 1776 838 1780
rect 930 1773 932 1777
rect 934 1773 936 1777
rect 948 1773 950 1777
rect 952 1773 954 1777
rect 967 1773 969 1777
rect 971 1773 973 1777
rect 527 1767 532 1771
rect 523 1764 532 1767
rect 535 1767 544 1771
rect 535 1764 548 1767
rect 556 1767 561 1771
rect 552 1764 561 1767
rect 563 1767 573 1771
rect 563 1764 577 1767
rect 585 1767 592 1771
rect 581 1764 592 1767
rect 595 1767 602 1771
rect 595 1764 606 1767
rect 614 1767 621 1771
rect 610 1764 621 1767
rect 624 1767 631 1771
rect 624 1764 635 1767
rect 643 1767 650 1771
rect 639 1764 650 1767
rect 653 1767 660 1771
rect 653 1764 664 1767
rect 672 1767 680 1771
rect 668 1764 680 1767
rect 683 1767 689 1771
rect 1381 1777 1385 1782
rect 1376 1773 1385 1777
rect 1389 1777 1395 1782
rect 1389 1773 1400 1777
rect 1412 1777 1417 1782
rect 1407 1773 1417 1777
rect 1421 1777 1426 1782
rect 1421 1773 1431 1777
rect 1445 1777 1451 1782
rect 1440 1773 1451 1777
rect 1455 1777 1459 1782
rect 1455 1773 1464 1777
rect 1556 1770 1558 1774
rect 1560 1770 1562 1774
rect 1574 1770 1576 1774
rect 1578 1770 1580 1774
rect 1593 1770 1595 1774
rect 1597 1770 1599 1774
rect 683 1764 693 1767
rect 1153 1764 1158 1768
rect 1149 1761 1158 1764
rect 1161 1764 1170 1768
rect 1161 1761 1174 1764
rect 1182 1764 1187 1768
rect 1178 1761 1187 1764
rect 1189 1764 1199 1768
rect 1189 1761 1203 1764
rect 1211 1764 1218 1768
rect 1207 1761 1218 1764
rect 1221 1764 1228 1768
rect 1221 1761 1232 1764
rect 1240 1764 1247 1768
rect 1236 1761 1247 1764
rect 1250 1764 1257 1768
rect 1250 1761 1261 1764
rect 1269 1764 1276 1768
rect 1265 1761 1276 1764
rect 1279 1764 1286 1768
rect 1279 1761 1290 1764
rect 1298 1764 1306 1768
rect 1294 1761 1306 1764
rect 1309 1764 1315 1768
rect 1981 1777 1985 1782
rect 1976 1773 1985 1777
rect 1989 1777 1995 1782
rect 1989 1773 2000 1777
rect 2012 1777 2017 1782
rect 2007 1773 2017 1777
rect 2021 1777 2026 1782
rect 2021 1773 2031 1777
rect 2045 1777 2051 1782
rect 2040 1773 2051 1777
rect 2055 1777 2059 1782
rect 2055 1773 2064 1777
rect 2156 1770 2158 1774
rect 2160 1770 2162 1774
rect 2174 1770 2176 1774
rect 2178 1770 2180 1774
rect 2193 1770 2195 1774
rect 2197 1770 2199 1774
rect 2584 1780 2588 1785
rect 2579 1776 2588 1780
rect 2592 1780 2598 1785
rect 2592 1776 2603 1780
rect 2615 1780 2620 1785
rect 2610 1776 2620 1780
rect 2624 1780 2629 1785
rect 2624 1776 2634 1780
rect 2648 1780 2654 1785
rect 2643 1776 2654 1780
rect 2658 1780 2662 1785
rect 2658 1776 2667 1780
rect 2759 1773 2761 1777
rect 2763 1773 2765 1777
rect 2777 1773 2779 1777
rect 2781 1773 2783 1777
rect 2796 1773 2798 1777
rect 2800 1773 2802 1777
rect 1309 1761 1319 1764
rect 1753 1764 1758 1768
rect 1749 1761 1758 1764
rect 1761 1764 1770 1768
rect 1761 1761 1774 1764
rect 1782 1764 1787 1768
rect 1778 1761 1787 1764
rect 1789 1764 1799 1768
rect 1789 1761 1803 1764
rect 1811 1764 1818 1768
rect 1807 1761 1818 1764
rect 1821 1764 1828 1768
rect 1821 1761 1832 1764
rect 1840 1764 1847 1768
rect 1836 1761 1847 1764
rect 1850 1764 1857 1768
rect 1850 1761 1861 1764
rect 1869 1764 1876 1768
rect 1865 1761 1876 1764
rect 1879 1764 1886 1768
rect 1879 1761 1890 1764
rect 1898 1764 1906 1768
rect 1894 1761 1906 1764
rect 1909 1764 1915 1768
rect 2356 1767 2361 1771
rect 2352 1764 2361 1767
rect 2364 1767 2373 1771
rect 2364 1764 2377 1767
rect 2385 1767 2390 1771
rect 2381 1764 2390 1767
rect 2392 1767 2402 1771
rect 2392 1764 2406 1767
rect 2414 1767 2421 1771
rect 2410 1765 2421 1767
rect 2413 1764 2421 1765
rect 2424 1767 2431 1771
rect 2424 1764 2435 1767
rect 2443 1767 2450 1771
rect 2439 1764 2450 1767
rect 2453 1767 2460 1771
rect 2453 1764 2464 1767
rect 2472 1767 2479 1771
rect 2468 1764 2479 1767
rect 2482 1767 2489 1771
rect 2482 1764 2493 1767
rect 2501 1767 2509 1771
rect 2497 1764 2509 1767
rect 2512 1767 2518 1771
rect 2512 1764 2522 1767
rect 1909 1761 1919 1764
rect 771 1641 775 1646
rect 766 1637 775 1641
rect 779 1641 785 1646
rect 779 1637 790 1641
rect 802 1641 807 1646
rect 797 1637 807 1641
rect 811 1641 816 1646
rect 811 1637 821 1641
rect 835 1641 841 1646
rect 830 1637 841 1641
rect 845 1641 849 1646
rect 845 1637 854 1641
rect 1397 1638 1401 1643
rect 1392 1634 1401 1638
rect 1405 1638 1411 1643
rect 1405 1634 1416 1638
rect 1428 1638 1433 1643
rect 1423 1634 1433 1638
rect 1437 1638 1442 1643
rect 1437 1634 1447 1638
rect 1461 1638 1467 1643
rect 1456 1634 1467 1638
rect 1471 1638 1475 1643
rect 1471 1634 1480 1638
rect 1997 1638 2001 1643
rect 1992 1634 2001 1638
rect 2005 1638 2011 1643
rect 2005 1634 2016 1638
rect 2028 1638 2033 1643
rect 2023 1634 2033 1638
rect 2037 1638 2042 1643
rect 2037 1634 2047 1638
rect 2061 1638 2067 1643
rect 2056 1634 2067 1638
rect 2071 1638 2075 1643
rect 2071 1634 2080 1638
rect 2600 1641 2604 1646
rect 2595 1637 2604 1641
rect 2608 1641 2614 1646
rect 2608 1637 2619 1641
rect 2631 1641 2636 1646
rect 2626 1637 2636 1641
rect 2640 1641 2645 1646
rect 2640 1637 2650 1641
rect 2664 1641 2670 1646
rect 2659 1637 2670 1641
rect 2674 1641 2678 1646
rect 2674 1637 2683 1641
rect 537 1511 542 1515
rect 533 1508 542 1511
rect 545 1511 554 1515
rect 545 1508 558 1511
rect 566 1511 571 1515
rect 562 1508 571 1511
rect 573 1511 583 1515
rect 573 1508 587 1511
rect 595 1511 602 1515
rect 591 1508 602 1511
rect 605 1511 612 1515
rect 605 1508 616 1511
rect 624 1511 631 1515
rect 620 1508 631 1511
rect 634 1511 641 1515
rect 634 1508 645 1511
rect 653 1511 660 1515
rect 649 1508 660 1511
rect 663 1511 670 1515
rect 663 1508 674 1511
rect 682 1511 690 1515
rect 678 1508 690 1511
rect 693 1511 699 1515
rect 693 1508 703 1511
rect 1163 1508 1168 1512
rect 1159 1505 1168 1508
rect 1171 1508 1180 1512
rect 1171 1505 1184 1508
rect 1192 1508 1197 1512
rect 1188 1505 1197 1508
rect 1199 1508 1209 1512
rect 1199 1505 1213 1508
rect 1221 1508 1228 1512
rect 1217 1505 1228 1508
rect 1231 1508 1238 1512
rect 1231 1505 1242 1508
rect 1250 1508 1257 1512
rect 1246 1505 1257 1508
rect 1260 1508 1267 1512
rect 1260 1505 1271 1508
rect 1279 1508 1286 1512
rect 1275 1505 1286 1508
rect 1289 1508 1296 1512
rect 1289 1505 1300 1508
rect 1308 1508 1316 1512
rect 1304 1505 1316 1508
rect 1319 1508 1325 1512
rect 1319 1505 1329 1508
rect 1763 1508 1768 1512
rect 1759 1505 1768 1508
rect 1771 1508 1780 1512
rect 1771 1505 1784 1508
rect 1792 1508 1797 1512
rect 1788 1505 1797 1508
rect 1799 1508 1809 1512
rect 1799 1505 1813 1508
rect 1821 1508 1828 1512
rect 1817 1505 1828 1508
rect 1831 1508 1838 1512
rect 1831 1505 1842 1508
rect 1850 1508 1857 1512
rect 1846 1505 1857 1508
rect 1860 1508 1867 1512
rect 1860 1505 1871 1508
rect 1879 1508 1886 1512
rect 1875 1505 1886 1508
rect 1889 1508 1896 1512
rect 1889 1505 1900 1508
rect 1908 1508 1916 1512
rect 1904 1505 1916 1508
rect 1919 1508 1925 1512
rect 2366 1511 2371 1515
rect 2362 1508 2371 1511
rect 2374 1511 2383 1515
rect 2374 1508 2387 1511
rect 2395 1511 2400 1515
rect 2391 1508 2400 1511
rect 2402 1511 2412 1515
rect 2402 1508 2416 1511
rect 2424 1511 2431 1515
rect 2420 1508 2431 1511
rect 2434 1511 2441 1515
rect 2434 1508 2445 1511
rect 2453 1511 2460 1515
rect 2449 1508 2460 1511
rect 2463 1511 2470 1515
rect 2463 1508 2474 1511
rect 2482 1511 2489 1515
rect 2478 1508 2489 1511
rect 2492 1511 2499 1515
rect 2492 1508 2503 1511
rect 2511 1511 2519 1515
rect 2507 1508 2519 1511
rect 2522 1511 2528 1515
rect 2522 1508 2532 1511
rect 1919 1505 1929 1508
rect 551 1150 556 1154
rect 547 1147 556 1150
rect 559 1150 568 1154
rect 559 1147 572 1150
rect 580 1150 585 1154
rect 576 1147 585 1150
rect 587 1150 597 1154
rect 587 1147 601 1150
rect 609 1150 616 1154
rect 605 1147 616 1150
rect 619 1150 626 1154
rect 619 1147 630 1150
rect 638 1150 645 1154
rect 634 1147 645 1150
rect 648 1150 655 1154
rect 648 1147 659 1150
rect 667 1150 674 1154
rect 663 1147 674 1150
rect 677 1150 684 1154
rect 677 1147 688 1150
rect 696 1150 704 1154
rect 692 1147 704 1150
rect 707 1150 713 1154
rect 707 1147 717 1150
rect 769 1150 774 1154
rect 765 1147 774 1150
rect 777 1150 786 1154
rect 777 1147 790 1150
rect 798 1150 803 1154
rect 794 1147 803 1150
rect 805 1150 815 1154
rect 805 1147 819 1150
rect 827 1150 834 1154
rect 823 1147 834 1150
rect 837 1150 844 1154
rect 837 1147 848 1150
rect 856 1150 863 1154
rect 852 1147 863 1150
rect 866 1150 873 1154
rect 866 1147 877 1150
rect 885 1150 892 1154
rect 881 1147 892 1150
rect 895 1150 902 1154
rect 895 1147 906 1150
rect 914 1150 922 1154
rect 910 1147 922 1150
rect 925 1150 931 1154
rect 925 1147 935 1150
rect 1002 1152 1007 1156
rect 998 1149 1007 1152
rect 1010 1152 1019 1156
rect 1010 1149 1023 1152
rect 1031 1152 1036 1156
rect 1027 1149 1036 1152
rect 1038 1152 1048 1156
rect 1038 1149 1052 1152
rect 1060 1152 1067 1156
rect 1056 1149 1067 1152
rect 1070 1152 1077 1156
rect 1070 1149 1081 1152
rect 1089 1152 1096 1156
rect 1085 1149 1096 1152
rect 1099 1152 1106 1156
rect 1099 1149 1110 1152
rect 1118 1152 1125 1156
rect 1114 1149 1125 1152
rect 1128 1152 1135 1156
rect 1128 1149 1139 1152
rect 1147 1152 1155 1156
rect 1143 1149 1155 1152
rect 1158 1152 1164 1156
rect 1158 1149 1168 1152
rect 1262 1153 1267 1157
rect 1258 1150 1267 1153
rect 1270 1153 1279 1157
rect 1270 1150 1283 1153
rect 1291 1153 1296 1157
rect 1287 1150 1296 1153
rect 1298 1153 1308 1157
rect 1298 1150 1312 1153
rect 1320 1153 1327 1157
rect 1316 1150 1327 1153
rect 1330 1153 1337 1157
rect 1330 1150 1341 1153
rect 1349 1153 1356 1157
rect 1345 1150 1356 1153
rect 1359 1153 1366 1157
rect 1359 1150 1370 1153
rect 1378 1153 1385 1157
rect 1374 1150 1385 1153
rect 1388 1153 1395 1157
rect 1388 1150 1399 1153
rect 1407 1153 1415 1157
rect 1403 1150 1415 1153
rect 1418 1153 1424 1157
rect 1418 1150 1428 1153
rect -405 1013 -401 1018
rect -410 1009 -401 1013
rect -397 1013 -391 1018
rect -397 1009 -386 1013
rect -374 1013 -369 1018
rect -379 1009 -369 1013
rect -365 1013 -360 1018
rect -365 1009 -355 1013
rect -341 1013 -335 1018
rect -346 1009 -335 1013
rect -331 1013 -327 1018
rect -331 1009 -322 1013
rect -269 1014 -265 1019
rect -274 1010 -265 1014
rect -261 1014 -255 1019
rect -261 1010 -250 1014
rect -238 1014 -233 1019
rect -243 1010 -233 1014
rect -229 1014 -224 1019
rect -229 1010 -219 1014
rect -205 1014 -199 1019
rect -210 1010 -199 1014
rect -195 1014 -191 1019
rect -195 1010 -186 1014
rect -134 1015 -130 1020
rect -139 1011 -130 1015
rect -126 1015 -120 1020
rect -126 1011 -115 1015
rect -103 1015 -98 1020
rect -108 1011 -98 1015
rect -94 1015 -89 1020
rect -94 1011 -84 1015
rect -70 1015 -64 1020
rect -75 1011 -64 1015
rect -60 1015 -56 1020
rect -60 1011 -51 1015
rect 3 1013 7 1018
rect -2 1009 7 1013
rect 11 1013 17 1018
rect 11 1009 22 1013
rect 34 1013 39 1018
rect 29 1009 39 1013
rect 43 1013 48 1018
rect 43 1009 53 1013
rect 67 1013 73 1018
rect 62 1009 73 1013
rect 77 1013 81 1018
rect 77 1009 86 1013
rect 808 965 812 970
rect 803 961 812 965
rect 816 965 822 970
rect 816 961 827 965
rect 839 965 844 970
rect 834 961 844 965
rect 848 965 853 970
rect 848 961 858 965
rect 872 965 878 970
rect 867 961 878 965
rect 882 965 886 970
rect 882 961 891 965
rect 983 958 985 962
rect 987 958 989 962
rect 1001 958 1003 962
rect 1005 958 1007 962
rect 1020 958 1022 962
rect 1024 958 1026 962
rect 580 952 585 956
rect -406 893 -402 898
rect -411 889 -402 893
rect -398 893 -392 898
rect -398 889 -387 893
rect -375 893 -370 898
rect -380 889 -370 893
rect -366 893 -361 898
rect -366 889 -356 893
rect -342 893 -336 898
rect -347 889 -336 893
rect -332 893 -328 898
rect -332 889 -323 893
rect -260 894 -256 899
rect -265 890 -256 894
rect -252 894 -246 899
rect -252 890 -241 894
rect -229 894 -224 899
rect -234 890 -224 894
rect -220 894 -215 899
rect -220 890 -210 894
rect -196 894 -190 899
rect -201 890 -190 894
rect -186 894 -182 899
rect -186 890 -177 894
rect -130 897 -126 902
rect -135 893 -126 897
rect -122 897 -116 902
rect -122 893 -111 897
rect -99 897 -94 902
rect -104 893 -94 897
rect -90 897 -85 902
rect -90 893 -80 897
rect -66 897 -60 902
rect -71 893 -60 897
rect -56 897 -52 902
rect 576 949 585 952
rect 588 952 597 956
rect 588 949 601 952
rect 609 952 614 956
rect 605 949 614 952
rect 616 952 626 956
rect 616 949 630 952
rect 638 952 645 956
rect 634 949 645 952
rect 648 952 655 956
rect 648 949 659 952
rect 667 952 674 956
rect 663 949 674 952
rect 677 952 684 956
rect 677 949 688 952
rect 696 952 703 956
rect 692 949 703 952
rect 706 952 713 956
rect 706 949 717 952
rect 725 952 733 956
rect 721 949 733 952
rect 736 952 742 956
rect 1434 962 1438 967
rect 1429 958 1438 962
rect 1442 962 1448 967
rect 1442 958 1453 962
rect 1465 962 1470 967
rect 1460 958 1470 962
rect 1474 962 1479 967
rect 1474 958 1484 962
rect 1498 962 1504 967
rect 1493 958 1504 962
rect 1508 962 1512 967
rect 1508 958 1517 962
rect 1609 955 1611 959
rect 1613 955 1615 959
rect 1627 955 1629 959
rect 1631 955 1633 959
rect 1646 955 1648 959
rect 1650 955 1652 959
rect 736 949 746 952
rect 1206 949 1211 953
rect 1202 946 1211 949
rect 1214 949 1223 953
rect 1214 946 1227 949
rect 1235 949 1240 953
rect 1231 946 1240 949
rect 1242 949 1252 953
rect 1242 946 1256 949
rect 1264 949 1271 953
rect 1260 946 1271 949
rect 1274 949 1281 953
rect 1274 946 1285 949
rect 1293 949 1300 953
rect 1289 946 1300 949
rect 1303 949 1310 953
rect 1303 946 1314 949
rect 1322 949 1329 953
rect 1318 946 1329 949
rect 1332 949 1339 953
rect 1332 946 1343 949
rect 1351 949 1359 953
rect 1347 946 1359 949
rect 1362 949 1368 953
rect 2034 962 2038 967
rect 2029 958 2038 962
rect 2042 962 2048 967
rect 2042 958 2053 962
rect 2065 962 2070 967
rect 2060 958 2070 962
rect 2074 962 2079 967
rect 2074 958 2084 962
rect 2098 962 2104 967
rect 2093 958 2104 962
rect 2108 962 2112 967
rect 2108 958 2117 962
rect 2209 955 2211 959
rect 2213 955 2215 959
rect 2227 955 2229 959
rect 2231 955 2233 959
rect 2246 955 2248 959
rect 2250 955 2252 959
rect 2637 965 2641 970
rect 2632 961 2641 965
rect 2645 965 2651 970
rect 2645 961 2656 965
rect 2668 965 2673 970
rect 2663 961 2673 965
rect 2677 965 2682 970
rect 2677 961 2687 965
rect 2701 965 2707 970
rect 2696 961 2707 965
rect 2711 965 2715 970
rect 2711 961 2720 965
rect 2812 958 2814 962
rect 2816 958 2818 962
rect 2830 958 2832 962
rect 2834 958 2836 962
rect 2849 958 2851 962
rect 2853 958 2855 962
rect 1362 946 1372 949
rect 1806 949 1811 953
rect 1802 946 1811 949
rect 1814 949 1823 953
rect 1814 946 1827 949
rect 1835 949 1840 953
rect 1831 946 1840 949
rect 1842 949 1852 953
rect 1842 946 1856 949
rect 1864 949 1871 953
rect 1860 946 1871 949
rect 1874 949 1881 953
rect 1874 946 1885 949
rect 1893 949 1900 953
rect 1889 946 1900 949
rect 1903 949 1910 953
rect 1903 946 1914 949
rect 1922 949 1929 953
rect 1918 946 1929 949
rect 1932 949 1939 953
rect 1932 946 1943 949
rect 1951 949 1959 953
rect 1947 946 1959 949
rect 1962 949 1968 953
rect 2409 952 2414 956
rect 2405 949 2414 952
rect 2417 952 2426 956
rect 2417 949 2430 952
rect 2438 952 2443 956
rect 2434 949 2443 952
rect 2445 952 2455 956
rect 2445 949 2459 952
rect 2467 952 2474 956
rect 2463 950 2474 952
rect 2466 949 2474 950
rect 2477 952 2484 956
rect 2477 949 2488 952
rect 2496 952 2503 956
rect 2492 949 2503 952
rect 2506 952 2513 956
rect 2506 949 2517 952
rect 2525 952 2532 956
rect 2521 949 2532 952
rect 2535 952 2542 956
rect 2535 949 2546 952
rect 2554 952 2562 956
rect 2550 949 2562 952
rect 2565 952 2571 956
rect 2565 949 2575 952
rect 1962 946 1972 949
rect -56 893 -47 897
rect 11 896 15 901
rect 6 892 15 896
rect 19 896 25 901
rect 19 892 30 896
rect 42 896 47 901
rect 37 892 47 896
rect 51 896 56 901
rect 51 892 61 896
rect 75 896 81 901
rect 70 892 81 896
rect 85 896 89 901
rect 85 892 94 896
rect 824 826 828 831
rect 819 822 828 826
rect 832 826 838 831
rect 832 822 843 826
rect 855 826 860 831
rect 850 822 860 826
rect 864 826 869 831
rect 864 822 874 826
rect 888 826 894 831
rect 883 822 894 826
rect 898 826 902 831
rect 898 822 907 826
rect 1450 823 1454 828
rect 1445 819 1454 823
rect 1458 823 1464 828
rect 1458 819 1469 823
rect 1481 823 1486 828
rect 1476 819 1486 823
rect 1490 823 1495 828
rect 1490 819 1500 823
rect 1514 823 1520 828
rect 1509 819 1520 823
rect 1524 823 1528 828
rect 1524 819 1533 823
rect 2050 823 2054 828
rect 2045 819 2054 823
rect 2058 823 2064 828
rect 2058 819 2069 823
rect 2081 823 2086 828
rect 2076 819 2086 823
rect 2090 823 2095 828
rect 2090 819 2100 823
rect 2114 823 2120 828
rect 2109 819 2120 823
rect 2124 823 2128 828
rect 2124 819 2133 823
rect 2653 826 2657 831
rect 2648 822 2657 826
rect 2661 826 2667 831
rect 2661 822 2672 826
rect 2684 826 2689 831
rect 2679 822 2689 826
rect 2693 826 2698 831
rect 2693 822 2703 826
rect 2717 826 2723 831
rect 2712 822 2723 826
rect 2727 826 2731 831
rect 2727 822 2736 826
rect 590 696 595 700
rect 586 693 595 696
rect 598 696 607 700
rect 598 693 611 696
rect 619 696 624 700
rect 615 693 624 696
rect 626 696 636 700
rect 626 693 640 696
rect 648 696 655 700
rect 644 693 655 696
rect 658 696 665 700
rect 658 693 669 696
rect 677 696 684 700
rect 673 693 684 696
rect 687 696 694 700
rect 687 693 698 696
rect 706 696 713 700
rect 702 693 713 696
rect 716 696 723 700
rect 716 693 727 696
rect 735 696 743 700
rect 731 693 743 696
rect 746 696 752 700
rect 746 693 756 696
rect 1216 693 1221 697
rect 1212 690 1221 693
rect 1224 693 1233 697
rect 1224 690 1237 693
rect 1245 693 1250 697
rect 1241 690 1250 693
rect 1252 693 1262 697
rect 1252 690 1266 693
rect 1274 693 1281 697
rect 1270 690 1281 693
rect 1284 693 1291 697
rect 1284 690 1295 693
rect 1303 693 1310 697
rect 1299 690 1310 693
rect 1313 693 1320 697
rect 1313 690 1324 693
rect 1332 693 1339 697
rect 1328 690 1339 693
rect 1342 693 1349 697
rect 1342 690 1353 693
rect 1361 693 1369 697
rect 1357 690 1369 693
rect 1372 693 1378 697
rect 1372 690 1382 693
rect 1816 693 1821 697
rect 1812 690 1821 693
rect 1824 693 1833 697
rect 1824 690 1837 693
rect 1845 693 1850 697
rect 1841 690 1850 693
rect 1852 693 1862 697
rect 1852 690 1866 693
rect 1874 693 1881 697
rect 1870 690 1881 693
rect 1884 693 1891 697
rect 1884 690 1895 693
rect 1903 693 1910 697
rect 1899 690 1910 693
rect 1913 693 1920 697
rect 1913 690 1924 693
rect 1932 693 1939 697
rect 1928 690 1939 693
rect 1942 693 1949 697
rect 1942 690 1953 693
rect 1961 693 1969 697
rect 1957 690 1969 693
rect 1972 693 1978 697
rect 2419 696 2424 700
rect 2415 693 2424 696
rect 2427 696 2436 700
rect 2427 693 2440 696
rect 2448 696 2453 700
rect 2444 693 2453 696
rect 2455 696 2465 700
rect 2455 693 2469 696
rect 2477 696 2484 700
rect 2473 693 2484 696
rect 2487 696 2494 700
rect 2487 693 2498 696
rect 2506 696 2513 700
rect 2502 693 2513 696
rect 2516 696 2523 700
rect 2516 693 2527 696
rect 2535 696 2542 700
rect 2531 693 2542 696
rect 2545 696 2552 700
rect 2545 693 2556 696
rect 2564 696 2572 700
rect 2560 693 2572 696
rect 2575 696 2581 700
rect 2575 693 2585 696
rect 1972 690 1982 693
rect -386 570 -382 575
rect -391 566 -382 570
rect -378 570 -372 575
rect -378 566 -367 570
rect -355 570 -350 575
rect -360 566 -350 570
rect -346 570 -341 575
rect -346 566 -336 570
rect -322 570 -316 575
rect -327 566 -316 570
rect -312 570 -308 575
rect -312 566 -303 570
rect -250 571 -246 576
rect -255 567 -246 571
rect -242 571 -236 576
rect -242 567 -231 571
rect -219 571 -214 576
rect -224 567 -214 571
rect -210 571 -205 576
rect -210 567 -200 571
rect -186 571 -180 576
rect -191 567 -180 571
rect -176 571 -172 576
rect -176 567 -167 571
rect -115 572 -111 577
rect -120 568 -111 572
rect -107 572 -101 577
rect -107 568 -96 572
rect -84 572 -79 577
rect -89 568 -79 572
rect -75 572 -70 577
rect -75 568 -65 572
rect -51 572 -45 577
rect -56 568 -45 572
rect -41 572 -37 577
rect -41 568 -32 572
rect 22 570 26 575
rect 17 566 26 570
rect 30 570 36 575
rect 30 566 41 570
rect 53 570 58 575
rect 48 566 58 570
rect 62 570 67 575
rect 62 566 72 570
rect 86 570 92 575
rect 81 566 92 570
rect 96 570 100 575
rect 96 566 105 570
rect -387 450 -383 455
rect -392 446 -383 450
rect -379 450 -373 455
rect -379 446 -368 450
rect -356 450 -351 455
rect -361 446 -351 450
rect -347 450 -342 455
rect -347 446 -337 450
rect -323 450 -317 455
rect -328 446 -317 450
rect -313 450 -309 455
rect -313 446 -304 450
rect -241 451 -237 456
rect -246 447 -237 451
rect -233 451 -227 456
rect -233 447 -222 451
rect -210 451 -205 456
rect -215 447 -205 451
rect -201 451 -196 456
rect -201 447 -191 451
rect -177 451 -171 456
rect -182 447 -171 451
rect -167 451 -163 456
rect -167 447 -158 451
rect -111 454 -107 459
rect -116 450 -107 454
rect -103 454 -97 459
rect -103 450 -92 454
rect -80 454 -75 459
rect -85 450 -75 454
rect -71 454 -66 459
rect -71 450 -61 454
rect -47 454 -41 459
rect -52 450 -41 454
rect -37 454 -33 459
rect -37 450 -28 454
rect 30 453 34 458
rect 25 449 34 453
rect 38 453 44 458
rect 38 449 49 453
rect 61 453 66 458
rect 56 449 66 453
rect 70 453 75 458
rect 70 449 80 453
rect 94 453 100 458
rect 89 449 100 453
rect 104 453 108 458
rect 104 449 113 453
rect -1047 396 -1043 401
rect -1052 392 -1043 396
rect -1039 396 -1033 401
rect -1039 392 -1028 396
rect -1016 396 -1011 401
rect -1021 392 -1011 396
rect -1007 396 -1002 401
rect -1007 392 -997 396
rect -983 396 -977 401
rect -988 392 -977 396
rect -973 396 -969 401
rect -973 392 -964 396
rect -1235 388 -1215 392
rect -1239 378 -1215 388
rect -1211 388 -1191 392
rect -1211 378 -1187 388
rect -1045 295 -1041 300
rect -1050 291 -1041 295
rect -1037 295 -1031 300
rect -1037 291 -1026 295
rect -1014 295 -1009 300
rect -1019 291 -1009 295
rect -1005 295 -1000 300
rect -1005 291 -995 295
rect -981 295 -975 300
rect -986 291 -975 295
rect -971 295 -967 300
rect -971 291 -962 295
rect -1042 196 -1038 201
rect -1047 192 -1038 196
rect -1034 196 -1028 201
rect -1034 192 -1023 196
rect -1011 196 -1006 201
rect -1016 192 -1006 196
rect -1002 196 -997 201
rect -1002 192 -992 196
rect -978 196 -972 201
rect -983 192 -972 196
rect -968 196 -964 201
rect -968 192 -959 196
rect -1237 169 -1217 173
rect -1241 159 -1217 169
rect -1213 169 -1193 173
rect -1213 159 -1189 169
rect -373 145 -369 150
rect -378 141 -369 145
rect -365 145 -359 150
rect -365 141 -354 145
rect -342 145 -337 150
rect -347 141 -337 145
rect -333 145 -328 150
rect -333 141 -323 145
rect -309 145 -303 150
rect -314 141 -303 145
rect -299 145 -295 150
rect -299 141 -290 145
rect -237 146 -233 151
rect -242 142 -233 146
rect -229 146 -223 151
rect -229 142 -218 146
rect -206 146 -201 151
rect -211 142 -201 146
rect -197 146 -192 151
rect -197 142 -187 146
rect -173 146 -167 151
rect -178 142 -167 146
rect -163 146 -159 151
rect -163 142 -154 146
rect -102 147 -98 152
rect -107 143 -98 147
rect -94 147 -88 152
rect -94 143 -83 147
rect -71 147 -66 152
rect -76 143 -66 147
rect -62 147 -57 152
rect -62 143 -52 147
rect -38 147 -32 152
rect -43 143 -32 147
rect -28 147 -24 152
rect -28 143 -19 147
rect 35 145 39 150
rect 30 141 39 145
rect 43 145 49 150
rect 43 141 54 145
rect 66 145 71 150
rect 61 141 71 145
rect 75 145 80 150
rect 75 141 85 145
rect 99 145 105 150
rect 94 141 105 145
rect 109 145 113 150
rect 109 141 118 145
rect -1040 88 -1036 93
rect -1045 84 -1036 88
rect -1032 88 -1026 93
rect -1032 84 -1021 88
rect -1009 88 -1004 93
rect -1014 84 -1004 88
rect -1000 88 -995 93
rect -1000 84 -990 88
rect -976 88 -970 93
rect -981 84 -970 88
rect -966 88 -962 93
rect -966 84 -957 88
rect -374 25 -370 30
rect -379 21 -370 25
rect -366 25 -360 30
rect -366 21 -355 25
rect -343 25 -338 30
rect -348 21 -338 25
rect -334 25 -329 30
rect -334 21 -324 25
rect -310 25 -304 30
rect -315 21 -304 25
rect -300 25 -296 30
rect -300 21 -291 25
rect -228 26 -224 31
rect -233 22 -224 26
rect -220 26 -214 31
rect -220 22 -209 26
rect -197 26 -192 31
rect -202 22 -192 26
rect -188 26 -183 31
rect -188 22 -178 26
rect -164 26 -158 31
rect -169 22 -158 26
rect -154 26 -150 31
rect -154 22 -145 26
rect -98 29 -94 34
rect -103 25 -94 29
rect -90 29 -84 34
rect -90 25 -79 29
rect -67 29 -62 34
rect -72 25 -62 29
rect -58 29 -53 34
rect -58 25 -48 29
rect -34 29 -28 34
rect -39 25 -28 29
rect -24 29 -20 34
rect -24 25 -15 29
rect 43 28 47 33
rect 38 24 47 28
rect 51 28 57 33
rect 51 24 62 28
rect 74 28 79 33
rect 69 24 79 28
rect 83 28 88 33
rect 83 24 93 28
rect 107 28 113 33
rect 102 24 113 28
rect 117 28 121 33
rect 117 24 126 28
rect 2081 -28 2101 -24
rect 2077 -38 2101 -28
rect 2105 -28 2125 -24
rect 2105 -38 2129 -28
rect 2606 -27 2626 -23
rect 2351 -33 2371 -29
rect 2347 -43 2371 -33
rect 2375 -33 2395 -29
rect 2375 -43 2399 -33
rect 2602 -37 2626 -27
rect 2630 -27 2650 -23
rect 2630 -37 2654 -27
rect 2874 -27 2894 -23
rect 2870 -37 2894 -27
rect 2898 -27 2918 -23
rect 2898 -37 2922 -27
rect -321 -305 -317 -300
rect -326 -309 -317 -305
rect -313 -305 -307 -300
rect -313 -309 -302 -305
rect -290 -305 -285 -300
rect -295 -309 -285 -305
rect -281 -305 -276 -300
rect -281 -309 -271 -305
rect -257 -305 -251 -300
rect -262 -309 -251 -305
rect -247 -305 -243 -300
rect -247 -309 -238 -305
rect -185 -304 -181 -299
rect -190 -308 -181 -304
rect -177 -304 -171 -299
rect -177 -308 -166 -304
rect -154 -304 -149 -299
rect -159 -308 -149 -304
rect -145 -304 -140 -299
rect -145 -308 -135 -304
rect -121 -304 -115 -299
rect -126 -308 -115 -304
rect -111 -304 -107 -299
rect -111 -308 -102 -304
rect -50 -303 -46 -298
rect -55 -307 -46 -303
rect -42 -303 -36 -298
rect -42 -307 -31 -303
rect -19 -303 -14 -298
rect -24 -307 -14 -303
rect -10 -303 -5 -298
rect -10 -307 0 -303
rect 14 -303 20 -298
rect 9 -307 20 -303
rect 24 -303 28 -298
rect 24 -307 33 -303
rect 87 -305 91 -300
rect 82 -309 91 -305
rect 95 -305 101 -300
rect 95 -309 106 -305
rect 118 -305 123 -300
rect 113 -309 123 -305
rect 127 -305 132 -300
rect 127 -309 137 -305
rect 151 -305 157 -300
rect 146 -309 157 -305
rect 161 -305 165 -300
rect 161 -309 170 -305
rect 3430 -219 3438 -215
rect 3426 -224 3438 -219
rect 3442 -219 3451 -215
rect 3442 -224 3455 -219
rect 3464 -219 3473 -215
rect 3460 -224 3473 -219
rect 3477 -219 3485 -215
rect 3477 -224 3489 -219
rect 3497 -219 3506 -215
rect 3493 -224 3506 -219
rect 3510 -219 3518 -215
rect 3510 -224 3522 -219
rect 3530 -219 3539 -215
rect 3526 -224 3539 -219
rect 3543 -219 3551 -215
rect 3543 -224 3555 -219
rect 3563 -219 3572 -215
rect 3559 -224 3572 -219
rect 3576 -219 3584 -215
rect 3576 -224 3588 -219
rect 2223 -290 2235 -286
rect 2219 -297 2235 -290
rect 2239 -290 2255 -286
rect 2239 -297 2259 -290
rect 2267 -290 2281 -286
rect 2263 -297 2281 -290
rect 2285 -290 2299 -286
rect 2285 -297 2303 -290
rect 2311 -290 2326 -286
rect 2307 -297 2326 -290
rect 2330 -290 2343 -286
rect 2330 -297 2347 -290
rect 2355 -290 2369 -286
rect 2351 -297 2369 -290
rect 2373 -290 2387 -286
rect 2373 -297 2391 -290
rect 2399 -290 2414 -286
rect 2395 -297 2414 -290
rect 2418 -290 2431 -286
rect 2418 -297 2435 -290
rect 2443 -290 2457 -286
rect 2439 -297 2457 -290
rect 2461 -290 2475 -286
rect 2461 -297 2479 -290
rect 2605 -290 2617 -286
rect 2601 -297 2617 -290
rect 2621 -290 2637 -286
rect 2621 -297 2641 -290
rect 2649 -290 2663 -286
rect 2645 -297 2663 -290
rect 2667 -290 2681 -286
rect 2667 -297 2685 -290
rect 2693 -290 2708 -286
rect 2689 -297 2708 -290
rect 2712 -290 2725 -286
rect 2712 -297 2729 -290
rect 2737 -290 2751 -286
rect 2733 -297 2751 -290
rect 2755 -290 2769 -286
rect 2755 -297 2773 -290
rect 2781 -290 2796 -286
rect 2777 -297 2796 -290
rect 2800 -290 2813 -286
rect 2800 -297 2817 -290
rect 2825 -290 2839 -286
rect 2821 -297 2839 -290
rect 2843 -290 2857 -286
rect 2843 -297 2861 -290
rect 2987 -290 2999 -286
rect 2983 -297 2999 -290
rect 3003 -290 3019 -286
rect 3003 -297 3023 -290
rect 3031 -290 3045 -286
rect 3027 -297 3045 -290
rect 3049 -290 3063 -286
rect 3049 -297 3067 -290
rect 3075 -290 3090 -286
rect 3071 -297 3090 -290
rect 3094 -290 3107 -286
rect 3094 -297 3111 -290
rect 3119 -290 3133 -286
rect 3115 -297 3133 -290
rect 3137 -290 3151 -286
rect 3137 -297 3155 -290
rect 3163 -290 3178 -286
rect 3159 -297 3178 -290
rect 3182 -290 3195 -286
rect 3182 -297 3199 -290
rect 3207 -290 3221 -286
rect 3203 -297 3221 -290
rect 3225 -290 3239 -286
rect 3225 -297 3243 -290
rect 2046 -317 2050 -312
rect 2041 -321 2050 -317
rect 2054 -317 2060 -312
rect 2054 -321 2065 -317
rect 2077 -317 2082 -312
rect 2072 -321 2082 -317
rect 2086 -317 2091 -312
rect 2086 -321 2096 -317
rect 2110 -317 2116 -312
rect 2105 -321 2116 -317
rect 2120 -317 2124 -312
rect 2120 -321 2129 -317
rect -322 -425 -318 -420
rect -327 -429 -318 -425
rect -314 -425 -308 -420
rect -314 -429 -303 -425
rect -291 -425 -286 -420
rect -296 -429 -286 -425
rect -282 -425 -277 -420
rect -282 -429 -272 -425
rect -258 -425 -252 -420
rect -263 -429 -252 -425
rect -248 -425 -244 -420
rect -248 -429 -239 -425
rect -176 -424 -172 -419
rect -181 -428 -172 -424
rect -168 -424 -162 -419
rect -168 -428 -157 -424
rect -145 -424 -140 -419
rect -150 -428 -140 -424
rect -136 -424 -131 -419
rect -136 -428 -126 -424
rect -112 -424 -106 -419
rect -117 -428 -106 -424
rect -102 -424 -98 -419
rect -102 -428 -93 -424
rect -46 -421 -42 -416
rect -51 -425 -42 -421
rect -38 -421 -32 -416
rect -38 -425 -27 -421
rect -15 -421 -10 -416
rect -20 -425 -10 -421
rect -6 -421 -1 -416
rect -6 -425 4 -421
rect 18 -421 24 -416
rect 13 -425 24 -421
rect 28 -421 32 -416
rect 28 -425 37 -421
rect 95 -422 99 -417
rect 90 -426 99 -422
rect 103 -422 109 -417
rect 103 -426 114 -422
rect 126 -422 131 -417
rect 121 -426 131 -422
rect 135 -422 140 -417
rect 135 -426 145 -422
rect 159 -422 165 -417
rect 154 -426 165 -422
rect 169 -422 173 -417
rect 169 -426 178 -422
rect 406 -485 410 -480
rect 401 -489 410 -485
rect 414 -485 420 -480
rect 414 -489 425 -485
rect 437 -485 442 -480
rect 432 -489 442 -485
rect 446 -485 451 -480
rect 446 -489 456 -485
rect 470 -485 476 -480
rect 465 -489 476 -485
rect 480 -485 484 -480
rect 480 -489 489 -485
rect -265 -591 -261 -586
rect -270 -595 -261 -591
rect -257 -591 -251 -586
rect -257 -595 -246 -591
rect -234 -591 -229 -586
rect -239 -595 -229 -591
rect -225 -591 -220 -586
rect -225 -595 -215 -591
rect -201 -591 -195 -586
rect -206 -595 -195 -591
rect -191 -591 -187 -586
rect -191 -595 -182 -591
rect 2061 -603 2067 -599
rect -89 -647 -85 -642
rect -94 -651 -85 -647
rect -81 -647 -75 -642
rect -81 -651 -70 -647
rect -58 -647 -53 -642
rect -63 -651 -53 -647
rect -49 -647 -44 -642
rect -49 -651 -39 -647
rect -25 -647 -19 -642
rect -30 -651 -19 -647
rect -15 -647 -11 -642
rect -15 -651 -6 -647
rect 2057 -605 2067 -603
rect 2070 -603 2080 -599
rect 2070 -605 2084 -603
rect 2095 -603 2102 -599
rect 2091 -605 2102 -603
rect 2105 -603 2114 -599
rect 2105 -605 2118 -603
rect 2128 -603 2137 -599
rect 2124 -605 2137 -603
rect 2140 -603 2147 -599
rect 2140 -605 2151 -603
rect 2160 -603 2169 -599
rect 2156 -605 2169 -603
rect 2172 -603 2179 -599
rect 2172 -605 2183 -603
rect 2192 -603 2200 -599
rect 2188 -605 2200 -603
rect 2203 -603 2211 -599
rect 2203 -605 2215 -603
rect 2224 -603 2233 -599
rect 2220 -605 2233 -603
rect 2236 -603 2243 -599
rect 2236 -605 2247 -603
rect 165 -657 169 -652
rect 160 -661 169 -657
rect 173 -657 179 -652
rect 173 -661 184 -657
rect 196 -657 201 -652
rect 191 -661 201 -657
rect 205 -657 210 -652
rect 205 -661 215 -657
rect 229 -657 235 -652
rect 224 -661 235 -657
rect 239 -657 243 -652
rect 239 -661 248 -657
rect 2060 -850 2066 -846
rect 2056 -852 2066 -850
rect 2069 -850 2079 -846
rect 2069 -852 2083 -850
rect 2094 -850 2101 -846
rect 2090 -852 2101 -850
rect 2104 -850 2113 -846
rect 2104 -852 2117 -850
rect 2127 -850 2136 -846
rect 2123 -852 2136 -850
rect 2139 -850 2146 -846
rect 2139 -852 2150 -850
rect 2159 -850 2168 -846
rect 2155 -852 2168 -850
rect 2171 -850 2178 -846
rect 2171 -852 2182 -850
rect 2191 -850 2199 -846
rect 2187 -852 2199 -850
rect 2202 -850 2210 -846
rect 2202 -852 2214 -850
rect 2223 -850 2232 -846
rect 2219 -852 2232 -850
rect 2235 -850 2242 -846
rect 2235 -852 2246 -850
rect 2414 -910 2426 -906
rect 2410 -917 2426 -910
rect 2430 -910 2446 -906
rect 2430 -917 2450 -910
rect 2458 -910 2472 -906
rect 2454 -917 2472 -910
rect 2476 -910 2490 -906
rect 2476 -917 2494 -910
rect 2502 -910 2517 -906
rect 2498 -917 2517 -910
rect 2521 -910 2534 -906
rect 2521 -917 2538 -910
rect 2546 -910 2560 -906
rect 2542 -917 2560 -910
rect 2564 -910 2578 -906
rect 2564 -917 2582 -910
rect 2590 -910 2605 -906
rect 2586 -917 2605 -910
rect 2609 -910 2622 -906
rect 2609 -917 2626 -910
rect 2634 -910 2648 -906
rect 2630 -917 2648 -910
rect 2652 -910 2666 -906
rect 2652 -917 2670 -910
rect 2064 -1076 2070 -1072
rect 2060 -1078 2070 -1076
rect 2073 -1076 2083 -1072
rect 2073 -1078 2087 -1076
rect 2098 -1076 2105 -1072
rect 2094 -1078 2105 -1076
rect 2108 -1076 2117 -1072
rect 2108 -1078 2121 -1076
rect 2131 -1076 2140 -1072
rect 2127 -1078 2140 -1076
rect 2143 -1076 2150 -1072
rect 2143 -1078 2154 -1076
rect 2163 -1076 2172 -1072
rect 2159 -1078 2172 -1076
rect 2175 -1076 2182 -1072
rect 2175 -1078 2186 -1076
rect 2195 -1076 2203 -1072
rect 2191 -1078 2203 -1076
rect 2206 -1076 2214 -1072
rect 2206 -1078 2218 -1076
rect 2227 -1076 2236 -1072
rect 2223 -1078 2236 -1076
rect 2239 -1076 2246 -1072
rect 2239 -1078 2250 -1076
rect 2061 -1283 2067 -1279
rect 2057 -1285 2067 -1283
rect 2070 -1283 2080 -1279
rect 2070 -1285 2084 -1283
rect 2095 -1283 2102 -1279
rect 2091 -1285 2102 -1283
rect 2105 -1283 2114 -1279
rect 2105 -1285 2118 -1283
rect 2128 -1283 2137 -1279
rect 2124 -1285 2137 -1283
rect 2140 -1283 2147 -1279
rect 2140 -1285 2151 -1283
rect 2160 -1283 2169 -1279
rect 2156 -1285 2169 -1283
rect 2172 -1283 2179 -1279
rect 2172 -1285 2183 -1283
rect 2192 -1283 2200 -1279
rect 2188 -1285 2200 -1283
rect 2203 -1283 2211 -1279
rect 2203 -1285 2215 -1283
rect 2224 -1283 2233 -1279
rect 2220 -1285 2233 -1283
rect 2236 -1283 2243 -1279
rect 2236 -1285 2247 -1283
rect 2089 -1462 2093 -1457
rect 2084 -1466 2093 -1462
rect 2097 -1462 2103 -1457
rect 2097 -1466 2108 -1462
rect 2120 -1462 2125 -1457
rect 2115 -1466 2125 -1462
rect 2129 -1462 2134 -1457
rect 2129 -1466 2139 -1462
rect 2153 -1462 2159 -1457
rect 2148 -1466 2159 -1462
rect 2163 -1462 2167 -1457
rect 2163 -1466 2172 -1462
rect 2274 -1516 2286 -1512
rect 2270 -1523 2286 -1516
rect 2290 -1516 2306 -1512
rect 2290 -1523 2310 -1516
rect 2318 -1516 2332 -1512
rect 2314 -1523 2332 -1516
rect 2336 -1516 2350 -1512
rect 2336 -1523 2354 -1516
rect 2362 -1516 2377 -1512
rect 2358 -1523 2377 -1516
rect 2381 -1516 2394 -1512
rect 2381 -1523 2398 -1516
rect 2406 -1516 2420 -1512
rect 2402 -1523 2420 -1516
rect 2424 -1516 2438 -1512
rect 2424 -1523 2442 -1516
rect 2450 -1516 2465 -1512
rect 2446 -1523 2465 -1516
rect 2469 -1516 2482 -1512
rect 2469 -1523 2486 -1516
rect 2494 -1516 2508 -1512
rect 2490 -1523 2508 -1516
rect 2512 -1516 2526 -1512
rect 2512 -1523 2530 -1516
rect 2646 -1515 2658 -1511
rect 2642 -1522 2658 -1515
rect 2662 -1515 2678 -1511
rect 2662 -1522 2682 -1515
rect 2690 -1515 2704 -1511
rect 2686 -1522 2704 -1515
rect 2708 -1515 2722 -1511
rect 2708 -1522 2726 -1515
rect 2734 -1515 2749 -1511
rect 2730 -1522 2749 -1515
rect 2753 -1515 2766 -1511
rect 2753 -1522 2770 -1515
rect 2778 -1515 2792 -1511
rect 2774 -1522 2792 -1515
rect 2796 -1515 2810 -1511
rect 2796 -1522 2814 -1515
rect 2822 -1515 2837 -1511
rect 2818 -1522 2837 -1515
rect 2841 -1515 2854 -1511
rect 2841 -1522 2858 -1515
rect 2866 -1515 2880 -1511
rect 2862 -1522 2880 -1515
rect 2884 -1515 2898 -1511
rect 2884 -1522 2902 -1515
rect 3020 -1515 3032 -1511
rect 3016 -1522 3032 -1515
rect 3036 -1515 3052 -1511
rect 3036 -1522 3056 -1515
rect 3064 -1515 3078 -1511
rect 3060 -1522 3078 -1515
rect 3082 -1515 3096 -1511
rect 3082 -1522 3100 -1515
rect 3108 -1515 3123 -1511
rect 3104 -1522 3123 -1515
rect 3127 -1515 3140 -1511
rect 3127 -1522 3144 -1515
rect 3152 -1515 3166 -1511
rect 3148 -1522 3166 -1515
rect 3170 -1515 3184 -1511
rect 3170 -1522 3188 -1515
rect 3196 -1515 3211 -1511
rect 3192 -1522 3211 -1515
rect 3215 -1515 3228 -1511
rect 3215 -1522 3232 -1515
rect 3240 -1515 3254 -1511
rect 3236 -1522 3254 -1515
rect 3258 -1515 3272 -1511
rect 3258 -1522 3276 -1515
rect 3480 -1546 3488 -1542
rect 3476 -1551 3488 -1546
rect 3492 -1546 3501 -1542
rect 3492 -1551 3505 -1546
rect 3514 -1546 3523 -1542
rect 3510 -1551 3523 -1546
rect 3527 -1546 3535 -1542
rect 3527 -1551 3539 -1546
rect 3547 -1546 3556 -1542
rect 3543 -1551 3556 -1546
rect 3560 -1546 3568 -1542
rect 3560 -1551 3572 -1546
rect 3580 -1546 3589 -1542
rect 3576 -1551 3589 -1546
rect 3593 -1546 3601 -1542
rect 3593 -1551 3605 -1546
rect 3613 -1546 3622 -1542
rect 3609 -1551 3622 -1546
rect 3626 -1546 3634 -1542
rect 3626 -1551 3638 -1546
rect 2108 -1567 2128 -1563
rect 2104 -1577 2128 -1567
rect 2132 -1567 2152 -1563
rect 2132 -1577 2156 -1567
rect 2305 -1613 2325 -1609
rect 2301 -1623 2325 -1613
rect 2329 -1613 2349 -1609
rect 2329 -1623 2353 -1613
rect 2713 -1637 2733 -1633
rect 2709 -1647 2733 -1637
rect 2737 -1637 2757 -1633
rect 2737 -1647 2761 -1637
rect 3140 -1636 3160 -1632
rect 3136 -1646 3160 -1636
rect 3164 -1636 3184 -1632
rect 3164 -1646 3188 -1636
<< pdiffusion >>
rect 498 2037 503 2041
rect 494 2034 503 2037
rect 506 2037 515 2041
rect 506 2034 519 2037
rect 527 2037 532 2041
rect 523 2034 532 2037
rect 534 2037 544 2041
rect 534 2034 548 2037
rect 556 2037 563 2041
rect 552 2034 563 2037
rect 566 2037 573 2041
rect 566 2034 577 2037
rect 585 2037 592 2041
rect 581 2034 592 2037
rect 595 2037 602 2041
rect 595 2034 606 2037
rect 614 2037 621 2041
rect 610 2034 621 2037
rect 624 2037 631 2041
rect 624 2034 635 2037
rect 643 2037 651 2041
rect 639 2034 651 2037
rect 654 2037 660 2041
rect 654 2034 664 2037
rect 716 2037 721 2041
rect 712 2034 721 2037
rect 724 2037 733 2041
rect 724 2034 737 2037
rect 745 2037 750 2041
rect 741 2034 750 2037
rect 752 2037 762 2041
rect 752 2034 766 2037
rect 774 2037 781 2041
rect 770 2034 781 2037
rect 784 2037 791 2041
rect 784 2034 795 2037
rect 803 2037 810 2041
rect 799 2034 810 2037
rect 813 2037 820 2041
rect 813 2034 824 2037
rect 832 2037 839 2041
rect 828 2034 839 2037
rect 842 2037 849 2041
rect 842 2034 853 2037
rect 861 2037 869 2041
rect 857 2034 869 2037
rect 872 2037 878 2041
rect 872 2034 882 2037
rect 949 2039 954 2043
rect 945 2036 954 2039
rect 957 2039 966 2043
rect 957 2036 970 2039
rect 978 2039 983 2043
rect 974 2036 983 2039
rect 985 2039 995 2043
rect 985 2036 999 2039
rect 1007 2039 1014 2043
rect 1003 2036 1014 2039
rect 1017 2039 1024 2043
rect 1017 2036 1028 2039
rect 1036 2039 1043 2043
rect 1032 2036 1043 2039
rect 1046 2039 1053 2043
rect 1046 2036 1057 2039
rect 1065 2039 1072 2043
rect 1061 2036 1072 2039
rect 1075 2039 1082 2043
rect 1075 2036 1086 2039
rect 1094 2039 1102 2043
rect 1090 2036 1102 2039
rect 1105 2039 1111 2043
rect 1105 2036 1115 2039
rect 1209 2040 1214 2044
rect 1205 2037 1214 2040
rect 1217 2040 1226 2044
rect 1217 2037 1230 2040
rect 1238 2040 1243 2044
rect 1234 2037 1243 2040
rect 1245 2040 1255 2044
rect 1245 2037 1259 2040
rect 1267 2040 1274 2044
rect 1263 2037 1274 2040
rect 1277 2040 1284 2044
rect 1277 2037 1288 2040
rect 1296 2040 1303 2044
rect 1292 2037 1303 2040
rect 1306 2040 1313 2044
rect 1306 2037 1317 2040
rect 1325 2040 1332 2044
rect 1321 2037 1332 2040
rect 1335 2040 1342 2044
rect 1335 2037 1346 2040
rect 1354 2040 1362 2044
rect 1350 2037 1362 2040
rect 1365 2040 1371 2044
rect 1365 2037 1375 2040
rect 527 1839 532 1843
rect 523 1836 532 1839
rect 535 1839 544 1843
rect 535 1836 548 1839
rect 556 1839 561 1843
rect 552 1836 561 1839
rect 563 1839 573 1843
rect 563 1836 577 1839
rect 585 1839 592 1843
rect 581 1836 592 1839
rect 595 1839 602 1843
rect 595 1836 606 1839
rect 614 1839 621 1843
rect 610 1836 621 1839
rect 624 1839 631 1843
rect 624 1836 635 1839
rect 643 1839 650 1843
rect 639 1836 650 1839
rect 653 1839 660 1843
rect 653 1836 664 1839
rect 672 1839 680 1843
rect 668 1836 680 1839
rect 683 1839 689 1843
rect 683 1836 693 1839
rect 755 1838 759 1843
rect 750 1834 759 1838
rect 763 1838 769 1843
rect 763 1834 774 1838
rect 786 1838 791 1843
rect 781 1834 791 1838
rect 795 1838 800 1843
rect 795 1834 805 1838
rect 819 1838 825 1843
rect 814 1834 825 1838
rect 829 1838 833 1843
rect 829 1834 838 1838
rect 1153 1836 1158 1840
rect 1149 1833 1158 1836
rect 1161 1836 1170 1840
rect 1161 1833 1174 1836
rect 1182 1836 1187 1840
rect 1178 1833 1187 1836
rect 1189 1836 1199 1840
rect 1189 1833 1203 1836
rect 1211 1836 1218 1840
rect 1207 1833 1218 1836
rect 1221 1836 1228 1840
rect 1221 1833 1232 1836
rect 1240 1836 1247 1840
rect 1236 1833 1247 1836
rect 1250 1836 1257 1840
rect 1250 1833 1261 1836
rect 1269 1836 1276 1840
rect 1265 1833 1276 1836
rect 1279 1836 1286 1840
rect 1279 1833 1290 1836
rect 1298 1836 1306 1840
rect 1294 1833 1306 1836
rect 1309 1836 1315 1840
rect 1309 1833 1319 1836
rect 1381 1835 1385 1840
rect 930 1814 932 1818
rect 934 1814 936 1818
rect 948 1814 950 1818
rect 952 1814 954 1818
rect 967 1814 969 1818
rect 971 1814 973 1818
rect 1376 1831 1385 1835
rect 1389 1835 1395 1840
rect 1389 1831 1400 1835
rect 1412 1835 1417 1840
rect 1407 1831 1417 1835
rect 1421 1835 1426 1840
rect 1421 1831 1431 1835
rect 1445 1835 1451 1840
rect 1440 1831 1451 1835
rect 1455 1835 1459 1840
rect 1455 1831 1464 1835
rect 1753 1836 1758 1840
rect 1749 1833 1758 1836
rect 1761 1836 1770 1840
rect 1761 1833 1774 1836
rect 1782 1836 1787 1840
rect 1778 1833 1787 1836
rect 1789 1836 1799 1840
rect 1789 1833 1803 1836
rect 1811 1836 1818 1840
rect 1807 1833 1818 1836
rect 1821 1836 1828 1840
rect 1821 1833 1832 1836
rect 1840 1836 1847 1840
rect 1836 1833 1847 1836
rect 1850 1836 1857 1840
rect 1850 1833 1861 1836
rect 1869 1836 1876 1840
rect 1865 1833 1876 1836
rect 1879 1836 1886 1840
rect 1879 1833 1890 1836
rect 1898 1836 1906 1840
rect 1894 1833 1906 1836
rect 1909 1836 1915 1840
rect 1909 1833 1919 1836
rect 1981 1835 1985 1840
rect 1556 1811 1558 1815
rect 1560 1811 1562 1815
rect 1574 1811 1576 1815
rect 1578 1811 1580 1815
rect 1593 1811 1595 1815
rect 1597 1811 1599 1815
rect 1976 1831 1985 1835
rect 1989 1835 1995 1840
rect 1989 1831 2000 1835
rect 2012 1835 2017 1840
rect 2007 1831 2017 1835
rect 2021 1835 2026 1840
rect 2021 1831 2031 1835
rect 2045 1835 2051 1840
rect 2040 1831 2051 1835
rect 2055 1835 2059 1840
rect 2356 1839 2361 1843
rect 2352 1836 2361 1839
rect 2364 1839 2373 1843
rect 2364 1836 2377 1839
rect 2385 1839 2390 1843
rect 2381 1836 2390 1839
rect 2392 1839 2402 1843
rect 2392 1836 2406 1839
rect 2414 1839 2421 1843
rect 2410 1836 2421 1839
rect 2424 1839 2431 1843
rect 2424 1836 2435 1839
rect 2443 1839 2450 1843
rect 2439 1836 2450 1839
rect 2453 1839 2460 1843
rect 2453 1836 2464 1839
rect 2472 1839 2479 1843
rect 2468 1836 2479 1839
rect 2482 1839 2489 1843
rect 2482 1836 2493 1839
rect 2501 1839 2509 1843
rect 2497 1836 2509 1839
rect 2512 1839 2518 1843
rect 2512 1836 2522 1839
rect 2584 1838 2588 1843
rect 2055 1831 2064 1835
rect 2156 1811 2158 1815
rect 2160 1811 2162 1815
rect 2174 1811 2176 1815
rect 2178 1811 2180 1815
rect 2193 1811 2195 1815
rect 2197 1811 2199 1815
rect 2579 1834 2588 1838
rect 2592 1838 2598 1843
rect 2592 1834 2603 1838
rect 2615 1838 2620 1843
rect 2610 1834 2620 1838
rect 2624 1838 2629 1843
rect 2624 1834 2634 1838
rect 2648 1838 2654 1843
rect 2643 1834 2654 1838
rect 2658 1838 2662 1843
rect 2658 1834 2667 1838
rect 2759 1814 2761 1818
rect 2763 1814 2765 1818
rect 2777 1814 2779 1818
rect 2781 1814 2783 1818
rect 2796 1814 2798 1818
rect 2800 1814 2802 1818
rect 771 1699 775 1704
rect 766 1695 775 1699
rect 779 1699 785 1704
rect 779 1695 790 1699
rect 802 1699 807 1704
rect 797 1695 807 1699
rect 811 1699 816 1704
rect 811 1695 821 1699
rect 835 1699 841 1704
rect 830 1695 841 1699
rect 845 1699 849 1704
rect 845 1695 854 1699
rect 1397 1696 1401 1701
rect 1392 1692 1401 1696
rect 1405 1696 1411 1701
rect 1405 1692 1416 1696
rect 1428 1696 1433 1701
rect 1423 1692 1433 1696
rect 1437 1696 1442 1701
rect 1437 1692 1447 1696
rect 1461 1696 1467 1701
rect 1456 1692 1467 1696
rect 1471 1696 1475 1701
rect 1471 1692 1480 1696
rect 1997 1696 2001 1701
rect 1992 1692 2001 1696
rect 2005 1696 2011 1701
rect 2005 1692 2016 1696
rect 2028 1696 2033 1701
rect 2023 1692 2033 1696
rect 2037 1696 2042 1701
rect 2037 1692 2047 1696
rect 2061 1696 2067 1701
rect 2056 1692 2067 1696
rect 2071 1696 2075 1701
rect 2071 1692 2080 1696
rect 2600 1699 2604 1704
rect 2595 1695 2604 1699
rect 2608 1699 2614 1704
rect 2608 1695 2619 1699
rect 2631 1699 2636 1704
rect 2626 1695 2636 1699
rect 2640 1699 2645 1704
rect 2640 1695 2650 1699
rect 2664 1699 2670 1704
rect 2659 1695 2670 1699
rect 2674 1699 2678 1704
rect 2674 1695 2683 1699
rect 537 1583 542 1587
rect 533 1580 542 1583
rect 545 1583 554 1587
rect 545 1580 558 1583
rect 566 1583 571 1587
rect 562 1580 571 1583
rect 573 1583 583 1587
rect 573 1580 587 1583
rect 595 1583 602 1587
rect 591 1580 602 1583
rect 605 1583 612 1587
rect 605 1580 616 1583
rect 624 1583 631 1587
rect 620 1580 631 1583
rect 634 1583 641 1587
rect 634 1580 645 1583
rect 653 1583 660 1587
rect 649 1580 660 1583
rect 663 1583 670 1587
rect 663 1580 674 1583
rect 682 1583 690 1587
rect 678 1580 690 1583
rect 693 1583 699 1587
rect 693 1580 703 1583
rect 1163 1580 1168 1584
rect 1159 1577 1168 1580
rect 1171 1580 1180 1584
rect 1171 1577 1184 1580
rect 1192 1580 1197 1584
rect 1188 1577 1197 1580
rect 1199 1580 1209 1584
rect 1199 1577 1213 1580
rect 1221 1580 1228 1584
rect 1217 1577 1228 1580
rect 1231 1580 1238 1584
rect 1231 1577 1242 1580
rect 1250 1580 1257 1584
rect 1246 1577 1257 1580
rect 1260 1580 1267 1584
rect 1260 1577 1271 1580
rect 1279 1580 1286 1584
rect 1275 1577 1286 1580
rect 1289 1580 1296 1584
rect 1289 1577 1300 1580
rect 1308 1580 1316 1584
rect 1304 1577 1316 1580
rect 1319 1580 1325 1584
rect 1319 1577 1329 1580
rect 1763 1580 1768 1584
rect 1759 1577 1768 1580
rect 1771 1580 1780 1584
rect 1771 1577 1784 1580
rect 1792 1580 1797 1584
rect 1788 1577 1797 1580
rect 1799 1580 1809 1584
rect 1799 1577 1813 1580
rect 1821 1580 1828 1584
rect 1817 1577 1828 1580
rect 1831 1580 1838 1584
rect 1831 1577 1842 1580
rect 1850 1580 1857 1584
rect 1846 1577 1857 1580
rect 1860 1580 1867 1584
rect 1860 1577 1871 1580
rect 1879 1580 1886 1584
rect 1875 1577 1886 1580
rect 1889 1580 1896 1584
rect 1889 1577 1900 1580
rect 1908 1580 1916 1584
rect 1904 1577 1916 1580
rect 1919 1580 1925 1584
rect 2366 1583 2371 1587
rect 2362 1580 2371 1583
rect 2374 1583 2383 1587
rect 2374 1580 2387 1583
rect 2395 1583 2400 1587
rect 2391 1580 2400 1583
rect 2402 1583 2412 1587
rect 2402 1580 2416 1583
rect 2424 1583 2431 1587
rect 2420 1580 2431 1583
rect 2434 1583 2441 1587
rect 2434 1580 2445 1583
rect 2453 1583 2460 1587
rect 2449 1580 2460 1583
rect 2463 1583 2470 1587
rect 2463 1580 2474 1583
rect 2482 1583 2489 1587
rect 2478 1580 2489 1583
rect 2492 1583 2499 1587
rect 2492 1580 2503 1583
rect 2511 1583 2519 1587
rect 2507 1580 2519 1583
rect 2522 1583 2528 1587
rect 2522 1580 2532 1583
rect 1919 1577 1929 1580
rect 551 1222 556 1226
rect 547 1219 556 1222
rect 559 1222 568 1226
rect 559 1219 572 1222
rect 580 1222 585 1226
rect 576 1219 585 1222
rect 587 1222 597 1226
rect 587 1219 601 1222
rect 609 1222 616 1226
rect 605 1219 616 1222
rect 619 1222 626 1226
rect 619 1219 630 1222
rect 638 1222 645 1226
rect 634 1219 645 1222
rect 648 1222 655 1226
rect 648 1219 659 1222
rect 667 1222 674 1226
rect 663 1219 674 1222
rect 677 1222 684 1226
rect 677 1219 688 1222
rect 696 1222 704 1226
rect 692 1219 704 1222
rect 707 1222 713 1226
rect 707 1219 717 1222
rect 769 1222 774 1226
rect 765 1219 774 1222
rect 777 1222 786 1226
rect 777 1219 790 1222
rect 798 1222 803 1226
rect 794 1219 803 1222
rect 805 1222 815 1226
rect 805 1219 819 1222
rect 827 1222 834 1226
rect 823 1219 834 1222
rect 837 1222 844 1226
rect 837 1219 848 1222
rect 856 1222 863 1226
rect 852 1219 863 1222
rect 866 1222 873 1226
rect 866 1219 877 1222
rect 885 1222 892 1226
rect 881 1219 892 1222
rect 895 1222 902 1226
rect 895 1219 906 1222
rect 914 1222 922 1226
rect 910 1219 922 1222
rect 925 1222 931 1226
rect 925 1219 935 1222
rect 1002 1224 1007 1228
rect 998 1221 1007 1224
rect 1010 1224 1019 1228
rect 1010 1221 1023 1224
rect 1031 1224 1036 1228
rect 1027 1221 1036 1224
rect 1038 1224 1048 1228
rect 1038 1221 1052 1224
rect 1060 1224 1067 1228
rect 1056 1221 1067 1224
rect 1070 1224 1077 1228
rect 1070 1221 1081 1224
rect 1089 1224 1096 1228
rect 1085 1221 1096 1224
rect 1099 1224 1106 1228
rect 1099 1221 1110 1224
rect 1118 1224 1125 1228
rect 1114 1221 1125 1224
rect 1128 1224 1135 1228
rect 1128 1221 1139 1224
rect 1147 1224 1155 1228
rect 1143 1221 1155 1224
rect 1158 1224 1164 1228
rect 1158 1221 1168 1224
rect 1262 1225 1267 1229
rect 1258 1222 1267 1225
rect 1270 1225 1279 1229
rect 1270 1222 1283 1225
rect 1291 1225 1296 1229
rect 1287 1222 1296 1225
rect 1298 1225 1308 1229
rect 1298 1222 1312 1225
rect 1320 1225 1327 1229
rect 1316 1222 1327 1225
rect 1330 1225 1337 1229
rect 1330 1222 1341 1225
rect 1349 1225 1356 1229
rect 1345 1222 1356 1225
rect 1359 1225 1366 1229
rect 1359 1222 1370 1225
rect 1378 1225 1385 1229
rect 1374 1222 1385 1225
rect 1388 1225 1395 1229
rect 1388 1222 1399 1225
rect 1407 1225 1415 1229
rect 1403 1222 1415 1225
rect 1418 1225 1424 1229
rect 1418 1222 1428 1225
rect -405 1071 -401 1076
rect -410 1067 -401 1071
rect -397 1071 -391 1076
rect -397 1067 -386 1071
rect -374 1071 -369 1076
rect -379 1067 -369 1071
rect -365 1071 -360 1076
rect -365 1067 -355 1071
rect -341 1071 -335 1076
rect -346 1067 -335 1071
rect -331 1071 -327 1076
rect -331 1067 -322 1071
rect -269 1072 -265 1077
rect -274 1068 -265 1072
rect -261 1072 -255 1077
rect -261 1068 -250 1072
rect -238 1072 -233 1077
rect -243 1068 -233 1072
rect -229 1072 -224 1077
rect -229 1068 -219 1072
rect -205 1072 -199 1077
rect -210 1068 -199 1072
rect -195 1072 -191 1077
rect -195 1068 -186 1072
rect -134 1073 -130 1078
rect -139 1069 -130 1073
rect -126 1073 -120 1078
rect -126 1069 -115 1073
rect -103 1073 -98 1078
rect -108 1069 -98 1073
rect -94 1073 -89 1078
rect -94 1069 -84 1073
rect -70 1073 -64 1078
rect -75 1069 -64 1073
rect -60 1073 -56 1078
rect -60 1069 -51 1073
rect 3 1071 7 1076
rect -2 1067 7 1071
rect 11 1071 17 1076
rect 11 1067 22 1071
rect 34 1071 39 1076
rect 29 1067 39 1071
rect 43 1071 48 1076
rect 43 1067 53 1071
rect 67 1071 73 1076
rect 62 1067 73 1071
rect 77 1071 81 1076
rect 77 1067 86 1071
rect 580 1024 585 1028
rect 576 1021 585 1024
rect 588 1024 597 1028
rect 588 1021 601 1024
rect 609 1024 614 1028
rect 605 1021 614 1024
rect 616 1024 626 1028
rect 616 1021 630 1024
rect 638 1024 645 1028
rect 634 1021 645 1024
rect 648 1024 655 1028
rect 648 1021 659 1024
rect 667 1024 674 1028
rect 663 1021 674 1024
rect 677 1024 684 1028
rect 677 1021 688 1024
rect 696 1024 703 1028
rect 692 1021 703 1024
rect 706 1024 713 1028
rect 706 1021 717 1024
rect 725 1024 733 1028
rect 721 1021 733 1024
rect 736 1024 742 1028
rect 736 1021 746 1024
rect 808 1023 812 1028
rect -406 951 -402 956
rect -411 947 -402 951
rect -398 951 -392 956
rect -398 947 -387 951
rect -375 951 -370 956
rect -380 947 -370 951
rect -366 951 -361 956
rect -366 947 -356 951
rect -342 951 -336 956
rect -347 947 -336 951
rect -332 951 -328 956
rect -332 947 -323 951
rect -260 952 -256 957
rect -265 948 -256 952
rect -252 952 -246 957
rect -252 948 -241 952
rect -229 952 -224 957
rect -234 948 -224 952
rect -220 952 -215 957
rect -220 948 -210 952
rect -196 952 -190 957
rect -201 948 -190 952
rect -186 952 -182 957
rect -186 948 -177 952
rect -130 955 -126 960
rect -135 951 -126 955
rect -122 955 -116 960
rect -122 951 -111 955
rect -99 955 -94 960
rect -104 951 -94 955
rect -90 955 -85 960
rect -90 951 -80 955
rect -66 955 -60 960
rect -71 951 -60 955
rect -56 955 -52 960
rect -56 951 -47 955
rect 11 954 15 959
rect 6 950 15 954
rect 19 954 25 959
rect 19 950 30 954
rect 42 954 47 959
rect 37 950 47 954
rect 51 954 56 959
rect 51 950 61 954
rect 75 954 81 959
rect 70 950 81 954
rect 85 954 89 959
rect 803 1019 812 1023
rect 816 1023 822 1028
rect 816 1019 827 1023
rect 839 1023 844 1028
rect 834 1019 844 1023
rect 848 1023 853 1028
rect 848 1019 858 1023
rect 872 1023 878 1028
rect 867 1019 878 1023
rect 882 1023 886 1028
rect 882 1019 891 1023
rect 1206 1021 1211 1025
rect 1202 1018 1211 1021
rect 1214 1021 1223 1025
rect 1214 1018 1227 1021
rect 1235 1021 1240 1025
rect 1231 1018 1240 1021
rect 1242 1021 1252 1025
rect 1242 1018 1256 1021
rect 1264 1021 1271 1025
rect 1260 1018 1271 1021
rect 1274 1021 1281 1025
rect 1274 1018 1285 1021
rect 1293 1021 1300 1025
rect 1289 1018 1300 1021
rect 1303 1021 1310 1025
rect 1303 1018 1314 1021
rect 1322 1021 1329 1025
rect 1318 1018 1329 1021
rect 1332 1021 1339 1025
rect 1332 1018 1343 1021
rect 1351 1021 1359 1025
rect 1347 1018 1359 1021
rect 1362 1021 1368 1025
rect 1362 1018 1372 1021
rect 1434 1020 1438 1025
rect 983 999 985 1003
rect 987 999 989 1003
rect 1001 999 1003 1003
rect 1005 999 1007 1003
rect 1020 999 1022 1003
rect 1024 999 1026 1003
rect 85 950 94 954
rect 1429 1016 1438 1020
rect 1442 1020 1448 1025
rect 1442 1016 1453 1020
rect 1465 1020 1470 1025
rect 1460 1016 1470 1020
rect 1474 1020 1479 1025
rect 1474 1016 1484 1020
rect 1498 1020 1504 1025
rect 1493 1016 1504 1020
rect 1508 1020 1512 1025
rect 1508 1016 1517 1020
rect 1806 1021 1811 1025
rect 1802 1018 1811 1021
rect 1814 1021 1823 1025
rect 1814 1018 1827 1021
rect 1835 1021 1840 1025
rect 1831 1018 1840 1021
rect 1842 1021 1852 1025
rect 1842 1018 1856 1021
rect 1864 1021 1871 1025
rect 1860 1018 1871 1021
rect 1874 1021 1881 1025
rect 1874 1018 1885 1021
rect 1893 1021 1900 1025
rect 1889 1018 1900 1021
rect 1903 1021 1910 1025
rect 1903 1018 1914 1021
rect 1922 1021 1929 1025
rect 1918 1018 1929 1021
rect 1932 1021 1939 1025
rect 1932 1018 1943 1021
rect 1951 1021 1959 1025
rect 1947 1018 1959 1021
rect 1962 1021 1968 1025
rect 1962 1018 1972 1021
rect 2034 1020 2038 1025
rect 1609 996 1611 1000
rect 1613 996 1615 1000
rect 1627 996 1629 1000
rect 1631 996 1633 1000
rect 1646 996 1648 1000
rect 1650 996 1652 1000
rect 2029 1016 2038 1020
rect 2042 1020 2048 1025
rect 2042 1016 2053 1020
rect 2065 1020 2070 1025
rect 2060 1016 2070 1020
rect 2074 1020 2079 1025
rect 2074 1016 2084 1020
rect 2098 1020 2104 1025
rect 2093 1016 2104 1020
rect 2108 1020 2112 1025
rect 2409 1024 2414 1028
rect 2405 1021 2414 1024
rect 2417 1024 2426 1028
rect 2417 1021 2430 1024
rect 2438 1024 2443 1028
rect 2434 1021 2443 1024
rect 2445 1024 2455 1028
rect 2445 1021 2459 1024
rect 2467 1024 2474 1028
rect 2463 1021 2474 1024
rect 2477 1024 2484 1028
rect 2477 1021 2488 1024
rect 2496 1024 2503 1028
rect 2492 1021 2503 1024
rect 2506 1024 2513 1028
rect 2506 1021 2517 1024
rect 2525 1024 2532 1028
rect 2521 1021 2532 1024
rect 2535 1024 2542 1028
rect 2535 1021 2546 1024
rect 2554 1024 2562 1028
rect 2550 1021 2562 1024
rect 2565 1024 2571 1028
rect 2565 1021 2575 1024
rect 2637 1023 2641 1028
rect 2108 1016 2117 1020
rect 2209 996 2211 1000
rect 2213 996 2215 1000
rect 2227 996 2229 1000
rect 2231 996 2233 1000
rect 2246 996 2248 1000
rect 2250 996 2252 1000
rect 2632 1019 2641 1023
rect 2645 1023 2651 1028
rect 2645 1019 2656 1023
rect 2668 1023 2673 1028
rect 2663 1019 2673 1023
rect 2677 1023 2682 1028
rect 2677 1019 2687 1023
rect 2701 1023 2707 1028
rect 2696 1019 2707 1023
rect 2711 1023 2715 1028
rect 2711 1019 2720 1023
rect 2812 999 2814 1003
rect 2816 999 2818 1003
rect 2830 999 2832 1003
rect 2834 999 2836 1003
rect 2849 999 2851 1003
rect 2853 999 2855 1003
rect 824 884 828 889
rect 819 880 828 884
rect 832 884 838 889
rect 832 880 843 884
rect 855 884 860 889
rect 850 880 860 884
rect 864 884 869 889
rect 864 880 874 884
rect 888 884 894 889
rect 883 880 894 884
rect 898 884 902 889
rect 898 880 907 884
rect 1450 881 1454 886
rect 1445 877 1454 881
rect 1458 881 1464 886
rect 1458 877 1469 881
rect 1481 881 1486 886
rect 1476 877 1486 881
rect 1490 881 1495 886
rect 1490 877 1500 881
rect 1514 881 1520 886
rect 1509 877 1520 881
rect 1524 881 1528 886
rect 1524 877 1533 881
rect 2050 881 2054 886
rect 2045 877 2054 881
rect 2058 881 2064 886
rect 2058 877 2069 881
rect 2081 881 2086 886
rect 2076 877 2086 881
rect 2090 881 2095 886
rect 2090 877 2100 881
rect 2114 881 2120 886
rect 2109 877 2120 881
rect 2124 881 2128 886
rect 2124 877 2133 881
rect 2653 884 2657 889
rect 2648 880 2657 884
rect 2661 884 2667 889
rect 2661 880 2672 884
rect 2684 884 2689 889
rect 2679 880 2689 884
rect 2693 884 2698 889
rect 2693 880 2703 884
rect 2717 884 2723 889
rect 2712 880 2723 884
rect 2727 884 2731 889
rect 2727 880 2736 884
rect 590 768 595 772
rect 586 765 595 768
rect 598 768 607 772
rect 598 765 611 768
rect 619 768 624 772
rect 615 765 624 768
rect 626 768 636 772
rect 626 765 640 768
rect 648 768 655 772
rect 644 765 655 768
rect 658 768 665 772
rect 658 765 669 768
rect 677 768 684 772
rect 673 765 684 768
rect 687 768 694 772
rect 687 765 698 768
rect 706 768 713 772
rect 702 765 713 768
rect 716 768 723 772
rect 716 765 727 768
rect 735 768 743 772
rect 731 765 743 768
rect 746 768 752 772
rect 746 765 756 768
rect 1216 765 1221 769
rect 1212 762 1221 765
rect 1224 765 1233 769
rect 1224 762 1237 765
rect 1245 765 1250 769
rect 1241 762 1250 765
rect 1252 765 1262 769
rect 1252 762 1266 765
rect 1274 765 1281 769
rect 1270 762 1281 765
rect 1284 765 1291 769
rect 1284 762 1295 765
rect 1303 765 1310 769
rect 1299 762 1310 765
rect 1313 765 1320 769
rect 1313 762 1324 765
rect 1332 765 1339 769
rect 1328 762 1339 765
rect 1342 765 1349 769
rect 1342 762 1353 765
rect 1361 765 1369 769
rect 1357 762 1369 765
rect 1372 765 1378 769
rect 1372 762 1382 765
rect 1816 765 1821 769
rect 1812 762 1821 765
rect 1824 765 1833 769
rect 1824 762 1837 765
rect 1845 765 1850 769
rect 1841 762 1850 765
rect 1852 765 1862 769
rect 1852 762 1866 765
rect 1874 765 1881 769
rect 1870 762 1881 765
rect 1884 765 1891 769
rect 1884 762 1895 765
rect 1903 765 1910 769
rect 1899 762 1910 765
rect 1913 765 1920 769
rect 1913 762 1924 765
rect 1932 765 1939 769
rect 1928 762 1939 765
rect 1942 765 1949 769
rect 1942 762 1953 765
rect 1961 765 1969 769
rect 1957 762 1969 765
rect 1972 765 1978 769
rect 2419 768 2424 772
rect 2415 765 2424 768
rect 2427 768 2436 772
rect 2427 765 2440 768
rect 2448 768 2453 772
rect 2444 765 2453 768
rect 2455 768 2465 772
rect 2455 765 2469 768
rect 2477 768 2484 772
rect 2473 765 2484 768
rect 2487 768 2494 772
rect 2487 765 2498 768
rect 2506 768 2513 772
rect 2502 765 2513 768
rect 2516 768 2523 772
rect 2516 765 2527 768
rect 2535 768 2542 772
rect 2531 765 2542 768
rect 2545 768 2552 772
rect 2545 765 2556 768
rect 2564 768 2572 772
rect 2560 765 2572 768
rect 2575 768 2581 772
rect 2575 765 2585 768
rect 1972 762 1982 765
rect -386 628 -382 633
rect -391 624 -382 628
rect -378 628 -372 633
rect -378 624 -367 628
rect -355 628 -350 633
rect -360 624 -350 628
rect -346 628 -341 633
rect -346 624 -336 628
rect -322 628 -316 633
rect -327 624 -316 628
rect -312 628 -308 633
rect -312 624 -303 628
rect -250 629 -246 634
rect -255 625 -246 629
rect -242 629 -236 634
rect -242 625 -231 629
rect -219 629 -214 634
rect -224 625 -214 629
rect -210 629 -205 634
rect -210 625 -200 629
rect -186 629 -180 634
rect -191 625 -180 629
rect -176 629 -172 634
rect -176 625 -167 629
rect -115 630 -111 635
rect -120 626 -111 630
rect -107 630 -101 635
rect -107 626 -96 630
rect -84 630 -79 635
rect -89 626 -79 630
rect -75 630 -70 635
rect -75 626 -65 630
rect -51 630 -45 635
rect -56 626 -45 630
rect -41 630 -37 635
rect -41 626 -32 630
rect 22 628 26 633
rect 17 624 26 628
rect 30 628 36 633
rect 30 624 41 628
rect 53 628 58 633
rect 48 624 58 628
rect 62 628 67 633
rect 62 624 72 628
rect 86 628 92 633
rect 81 624 92 628
rect 96 628 100 633
rect 96 624 105 628
rect -387 508 -383 513
rect -392 504 -383 508
rect -379 508 -373 513
rect -379 504 -368 508
rect -356 508 -351 513
rect -361 504 -351 508
rect -347 508 -342 513
rect -347 504 -337 508
rect -323 508 -317 513
rect -328 504 -317 508
rect -313 508 -309 513
rect -313 504 -304 508
rect -241 509 -237 514
rect -246 505 -237 509
rect -233 509 -227 514
rect -233 505 -222 509
rect -210 509 -205 514
rect -215 505 -205 509
rect -201 509 -196 514
rect -201 505 -191 509
rect -177 509 -171 514
rect -182 505 -171 509
rect -167 509 -163 514
rect -167 505 -158 509
rect -111 512 -107 517
rect -116 508 -107 512
rect -103 512 -97 517
rect -103 508 -92 512
rect -80 512 -75 517
rect -85 508 -75 512
rect -71 512 -66 517
rect -71 508 -61 512
rect -47 512 -41 517
rect -52 508 -41 512
rect -37 512 -33 517
rect -37 508 -28 512
rect 30 511 34 516
rect -1047 454 -1043 459
rect -1052 450 -1043 454
rect -1039 454 -1033 459
rect -1039 450 -1028 454
rect -1016 454 -1011 459
rect -1021 450 -1011 454
rect -1007 454 -1002 459
rect -1007 450 -997 454
rect -983 454 -977 459
rect -988 450 -977 454
rect -973 454 -969 459
rect 25 507 34 511
rect 38 511 44 516
rect 38 507 49 511
rect 61 511 66 516
rect 56 507 66 511
rect 70 511 75 516
rect 70 507 80 511
rect 94 511 100 516
rect 89 507 100 511
rect 104 511 108 516
rect 104 507 113 511
rect -973 450 -964 454
rect -1235 426 -1215 430
rect -1239 420 -1215 426
rect -1211 426 -1191 430
rect -1211 420 -1187 426
rect -1045 353 -1041 358
rect -1050 349 -1041 353
rect -1037 353 -1031 358
rect -1037 349 -1026 353
rect -1014 353 -1009 358
rect -1019 349 -1009 353
rect -1005 353 -1000 358
rect -1005 349 -995 353
rect -981 353 -975 358
rect -986 349 -975 353
rect -971 353 -967 358
rect -971 349 -962 353
rect -1042 254 -1038 259
rect -1047 250 -1038 254
rect -1034 254 -1028 259
rect -1034 250 -1023 254
rect -1011 254 -1006 259
rect -1016 250 -1006 254
rect -1002 254 -997 259
rect -1002 250 -992 254
rect -978 254 -972 259
rect -983 250 -972 254
rect -968 254 -964 259
rect -968 250 -959 254
rect -1237 207 -1217 211
rect -1241 201 -1217 207
rect -1213 207 -1193 211
rect -1213 201 -1189 207
rect -373 203 -369 208
rect -378 199 -369 203
rect -365 203 -359 208
rect -365 199 -354 203
rect -342 203 -337 208
rect -347 199 -337 203
rect -333 203 -328 208
rect -333 199 -323 203
rect -309 203 -303 208
rect -314 199 -303 203
rect -299 203 -295 208
rect -299 199 -290 203
rect -237 204 -233 209
rect -242 200 -233 204
rect -229 204 -223 209
rect -229 200 -218 204
rect -206 204 -201 209
rect -211 200 -201 204
rect -197 204 -192 209
rect -197 200 -187 204
rect -173 204 -167 209
rect -178 200 -167 204
rect -163 204 -159 209
rect -163 200 -154 204
rect -102 205 -98 210
rect -107 201 -98 205
rect -94 205 -88 210
rect -94 201 -83 205
rect -71 205 -66 210
rect -76 201 -66 205
rect -62 205 -57 210
rect -62 201 -52 205
rect -38 205 -32 210
rect -43 201 -32 205
rect -28 205 -24 210
rect -28 201 -19 205
rect 35 203 39 208
rect -1040 146 -1036 151
rect -1045 142 -1036 146
rect -1032 146 -1026 151
rect -1032 142 -1021 146
rect -1009 146 -1004 151
rect -1014 142 -1004 146
rect -1000 146 -995 151
rect -1000 142 -990 146
rect -976 146 -970 151
rect -981 142 -970 146
rect -966 146 -962 151
rect 30 199 39 203
rect 43 203 49 208
rect 43 199 54 203
rect 66 203 71 208
rect 61 199 71 203
rect 75 203 80 208
rect 75 199 85 203
rect 99 203 105 208
rect 94 199 105 203
rect 109 203 113 208
rect 109 199 118 203
rect -966 142 -957 146
rect -374 83 -370 88
rect -379 79 -370 83
rect -366 83 -360 88
rect -366 79 -355 83
rect -343 83 -338 88
rect -348 79 -338 83
rect -334 83 -329 88
rect -334 79 -324 83
rect -310 83 -304 88
rect -315 79 -304 83
rect -300 83 -296 88
rect -300 79 -291 83
rect -228 84 -224 89
rect -233 80 -224 84
rect -220 84 -214 89
rect -220 80 -209 84
rect -197 84 -192 89
rect -202 80 -192 84
rect -188 84 -183 89
rect -188 80 -178 84
rect -164 84 -158 89
rect -169 80 -158 84
rect -154 84 -150 89
rect -154 80 -145 84
rect -98 87 -94 92
rect -103 83 -94 87
rect -90 87 -84 92
rect -90 83 -79 87
rect -67 87 -62 92
rect -72 83 -62 87
rect -58 87 -53 92
rect -58 83 -48 87
rect -34 87 -28 92
rect -39 83 -28 87
rect -24 87 -20 92
rect -24 83 -15 87
rect 43 86 47 91
rect 38 82 47 86
rect 51 86 57 91
rect 51 82 62 86
rect 74 86 79 91
rect 69 82 79 86
rect 83 86 88 91
rect 83 82 93 86
rect 107 86 113 91
rect 102 82 113 86
rect 117 86 121 91
rect 117 82 126 86
rect 2081 10 2101 14
rect 2077 4 2101 10
rect 2105 10 2125 14
rect 2105 4 2129 10
rect 2606 11 2626 15
rect 2351 5 2371 9
rect 2347 -1 2371 5
rect 2375 5 2395 9
rect 2602 5 2626 11
rect 2630 11 2650 15
rect 2630 5 2654 11
rect 2874 11 2894 15
rect 2870 5 2894 11
rect 2898 11 2918 15
rect 2898 5 2922 11
rect 2375 -1 2399 5
rect 3430 -137 3438 -133
rect 3426 -142 3438 -137
rect 3442 -137 3451 -133
rect 3442 -142 3455 -137
rect 3464 -137 3473 -133
rect 3460 -142 3473 -137
rect 3477 -137 3485 -133
rect 3477 -142 3489 -137
rect 3497 -137 3506 -133
rect 3493 -142 3506 -137
rect 3510 -137 3518 -133
rect 3510 -142 3522 -137
rect 3530 -137 3539 -133
rect 3526 -142 3539 -137
rect 3543 -137 3551 -133
rect 3543 -142 3555 -137
rect 3563 -137 3572 -133
rect 3559 -142 3572 -137
rect 3576 -137 3584 -133
rect 3576 -142 3588 -137
rect 2223 -187 2235 -183
rect 2219 -194 2235 -187
rect 2239 -187 2255 -183
rect 2239 -194 2259 -187
rect 2267 -187 2281 -183
rect 2263 -194 2281 -187
rect 2285 -187 2299 -183
rect 2285 -194 2303 -187
rect 2311 -187 2326 -183
rect 2307 -194 2326 -187
rect 2330 -187 2343 -183
rect 2330 -194 2347 -187
rect 2355 -187 2369 -183
rect 2351 -194 2369 -187
rect 2373 -187 2387 -183
rect 2373 -194 2391 -187
rect 2399 -187 2414 -183
rect 2395 -194 2414 -187
rect 2418 -187 2431 -183
rect 2418 -194 2435 -187
rect 2443 -187 2457 -183
rect 2439 -194 2457 -187
rect 2461 -187 2475 -183
rect 2461 -194 2479 -187
rect 2605 -187 2617 -183
rect 2601 -194 2617 -187
rect 2621 -187 2637 -183
rect 2621 -194 2641 -187
rect 2649 -187 2663 -183
rect 2645 -194 2663 -187
rect 2667 -187 2681 -183
rect 2667 -194 2685 -187
rect 2693 -187 2708 -183
rect 2689 -194 2708 -187
rect 2712 -187 2725 -183
rect 2712 -194 2729 -187
rect 2737 -187 2751 -183
rect 2733 -194 2751 -187
rect 2755 -187 2769 -183
rect 2755 -194 2773 -187
rect 2781 -187 2796 -183
rect 2777 -194 2796 -187
rect 2800 -187 2813 -183
rect 2800 -194 2817 -187
rect 2825 -187 2839 -183
rect 2821 -194 2839 -187
rect 2843 -187 2857 -183
rect 2843 -194 2861 -187
rect 2987 -187 2999 -183
rect 2983 -194 2999 -187
rect 3003 -187 3019 -183
rect 3003 -194 3023 -187
rect 3031 -187 3045 -183
rect 3027 -194 3045 -187
rect 3049 -187 3063 -183
rect 3049 -194 3067 -187
rect 3075 -187 3090 -183
rect 3071 -194 3090 -187
rect 3094 -187 3107 -183
rect 3094 -194 3111 -187
rect 3119 -187 3133 -183
rect 3115 -194 3133 -187
rect 3137 -187 3151 -183
rect 3137 -194 3155 -187
rect 3163 -187 3178 -183
rect 3159 -194 3178 -187
rect 3182 -187 3195 -183
rect 3182 -194 3199 -187
rect 3207 -187 3221 -183
rect 3203 -194 3221 -187
rect 3225 -187 3239 -183
rect 3225 -194 3243 -187
rect -321 -247 -317 -242
rect -326 -251 -317 -247
rect -313 -247 -307 -242
rect -313 -251 -302 -247
rect -290 -247 -285 -242
rect -295 -251 -285 -247
rect -281 -247 -276 -242
rect -281 -251 -271 -247
rect -257 -247 -251 -242
rect -262 -251 -251 -247
rect -247 -247 -243 -242
rect -247 -251 -238 -247
rect -185 -246 -181 -241
rect -190 -250 -181 -246
rect -177 -246 -171 -241
rect -177 -250 -166 -246
rect -154 -246 -149 -241
rect -159 -250 -149 -246
rect -145 -246 -140 -241
rect -145 -250 -135 -246
rect -121 -246 -115 -241
rect -126 -250 -115 -246
rect -111 -246 -107 -241
rect -111 -250 -102 -246
rect -50 -245 -46 -240
rect -55 -249 -46 -245
rect -42 -245 -36 -240
rect -42 -249 -31 -245
rect -19 -245 -14 -240
rect -24 -249 -14 -245
rect -10 -245 -5 -240
rect -10 -249 0 -245
rect 14 -245 20 -240
rect 9 -249 20 -245
rect 24 -245 28 -240
rect 24 -249 33 -245
rect 87 -247 91 -242
rect 82 -251 91 -247
rect 95 -247 101 -242
rect 95 -251 106 -247
rect 118 -247 123 -242
rect 113 -251 123 -247
rect 127 -247 132 -242
rect 127 -251 137 -247
rect 151 -247 157 -242
rect 146 -251 157 -247
rect 161 -247 165 -242
rect 161 -251 170 -247
rect 2046 -259 2050 -254
rect 2041 -263 2050 -259
rect 2054 -259 2060 -254
rect 2054 -263 2065 -259
rect 2077 -259 2082 -254
rect 2072 -263 2082 -259
rect 2086 -259 2091 -254
rect 2086 -263 2096 -259
rect 2110 -259 2116 -254
rect 2105 -263 2116 -259
rect 2120 -259 2124 -254
rect 2120 -263 2129 -259
rect -322 -367 -318 -362
rect -327 -371 -318 -367
rect -314 -367 -308 -362
rect -314 -371 -303 -367
rect -291 -367 -286 -362
rect -296 -371 -286 -367
rect -282 -367 -277 -362
rect -282 -371 -272 -367
rect -258 -367 -252 -362
rect -263 -371 -252 -367
rect -248 -367 -244 -362
rect -248 -371 -239 -367
rect -176 -366 -172 -361
rect -181 -370 -172 -366
rect -168 -366 -162 -361
rect -168 -370 -157 -366
rect -145 -366 -140 -361
rect -150 -370 -140 -366
rect -136 -366 -131 -361
rect -136 -370 -126 -366
rect -112 -366 -106 -361
rect -117 -370 -106 -366
rect -102 -366 -98 -361
rect -102 -370 -93 -366
rect -46 -363 -42 -358
rect -51 -367 -42 -363
rect -38 -363 -32 -358
rect -38 -367 -27 -363
rect -15 -363 -10 -358
rect -20 -367 -10 -363
rect -6 -363 -1 -358
rect -6 -367 4 -363
rect 18 -363 24 -358
rect 13 -367 24 -363
rect 28 -363 32 -358
rect 28 -367 37 -363
rect 95 -364 99 -359
rect 90 -368 99 -364
rect 103 -364 109 -359
rect 103 -368 114 -364
rect 126 -364 131 -359
rect 121 -368 131 -364
rect 135 -364 140 -359
rect 135 -368 145 -364
rect 159 -364 165 -359
rect 154 -368 165 -364
rect 169 -364 173 -359
rect 169 -368 178 -364
rect 406 -427 410 -422
rect 401 -431 410 -427
rect 414 -427 420 -422
rect 414 -431 425 -427
rect 437 -427 442 -422
rect 432 -431 442 -427
rect 446 -427 451 -422
rect 446 -431 456 -427
rect 470 -427 476 -422
rect 465 -431 476 -427
rect 480 -427 484 -422
rect 480 -431 489 -427
rect 2061 -514 2067 -510
rect 2057 -516 2067 -514
rect 2070 -514 2080 -510
rect 2070 -516 2084 -514
rect 2095 -514 2102 -510
rect 2091 -516 2102 -514
rect 2105 -514 2114 -510
rect 2105 -516 2118 -514
rect 2128 -514 2137 -510
rect 2124 -516 2137 -514
rect 2140 -514 2147 -510
rect 2140 -516 2151 -514
rect 2160 -514 2169 -510
rect 2156 -516 2169 -514
rect 2172 -514 2179 -510
rect 2172 -516 2183 -514
rect 2192 -514 2200 -510
rect 2188 -516 2200 -514
rect 2203 -514 2211 -510
rect 2203 -516 2215 -514
rect 2224 -514 2233 -510
rect 2220 -516 2233 -514
rect 2236 -514 2243 -510
rect 2236 -516 2247 -514
rect -265 -533 -261 -528
rect -270 -537 -261 -533
rect -257 -533 -251 -528
rect -257 -537 -246 -533
rect -234 -533 -229 -528
rect -239 -537 -229 -533
rect -225 -533 -220 -528
rect -225 -537 -215 -533
rect -201 -533 -195 -528
rect -206 -537 -195 -533
rect -191 -533 -187 -528
rect -191 -537 -182 -533
rect -89 -589 -85 -584
rect -94 -593 -85 -589
rect -81 -589 -75 -584
rect -81 -593 -70 -589
rect -58 -589 -53 -584
rect -63 -593 -53 -589
rect -49 -589 -44 -584
rect -49 -593 -39 -589
rect -25 -589 -19 -584
rect -30 -593 -19 -589
rect -15 -589 -11 -584
rect -15 -593 -6 -589
rect 165 -599 169 -594
rect 160 -603 169 -599
rect 173 -599 179 -594
rect 173 -603 184 -599
rect 196 -599 201 -594
rect 191 -603 201 -599
rect 205 -599 210 -594
rect 205 -603 215 -599
rect 229 -599 235 -594
rect 224 -603 235 -599
rect 239 -599 243 -594
rect 239 -603 248 -599
rect 2060 -761 2066 -757
rect 2056 -763 2066 -761
rect 2069 -761 2079 -757
rect 2069 -763 2083 -761
rect 2094 -761 2101 -757
rect 2090 -763 2101 -761
rect 2104 -761 2113 -757
rect 2104 -763 2117 -761
rect 2127 -761 2136 -757
rect 2123 -763 2136 -761
rect 2139 -761 2146 -757
rect 2139 -763 2150 -761
rect 2159 -761 2168 -757
rect 2155 -763 2168 -761
rect 2171 -761 2178 -757
rect 2171 -763 2182 -761
rect 2191 -761 2199 -757
rect 2187 -763 2199 -761
rect 2202 -761 2210 -757
rect 2202 -763 2214 -761
rect 2223 -761 2232 -757
rect 2219 -763 2232 -761
rect 2235 -761 2242 -757
rect 2235 -763 2246 -761
rect 2414 -807 2426 -803
rect 2410 -814 2426 -807
rect 2430 -807 2446 -803
rect 2430 -814 2450 -807
rect 2458 -807 2472 -803
rect 2454 -814 2472 -807
rect 2476 -807 2490 -803
rect 2476 -814 2494 -807
rect 2502 -807 2517 -803
rect 2498 -814 2517 -807
rect 2521 -807 2534 -803
rect 2521 -814 2538 -807
rect 2546 -807 2560 -803
rect 2542 -814 2560 -807
rect 2564 -807 2578 -803
rect 2564 -814 2582 -807
rect 2590 -807 2605 -803
rect 2586 -814 2605 -807
rect 2609 -807 2622 -803
rect 2609 -814 2626 -807
rect 2634 -807 2648 -803
rect 2630 -814 2648 -807
rect 2652 -807 2666 -803
rect 2652 -814 2670 -807
rect 2064 -987 2070 -983
rect 2060 -989 2070 -987
rect 2073 -987 2083 -983
rect 2073 -989 2087 -987
rect 2098 -987 2105 -983
rect 2094 -989 2105 -987
rect 2108 -987 2117 -983
rect 2108 -989 2121 -987
rect 2131 -987 2140 -983
rect 2127 -989 2140 -987
rect 2143 -987 2150 -983
rect 2143 -989 2154 -987
rect 2163 -987 2172 -983
rect 2159 -989 2172 -987
rect 2175 -987 2182 -983
rect 2175 -989 2186 -987
rect 2195 -987 2203 -983
rect 2191 -989 2203 -987
rect 2206 -987 2214 -983
rect 2206 -989 2218 -987
rect 2227 -987 2236 -983
rect 2223 -989 2236 -987
rect 2239 -987 2246 -983
rect 2239 -989 2250 -987
rect 2061 -1194 2067 -1190
rect 2057 -1196 2067 -1194
rect 2070 -1194 2080 -1190
rect 2070 -1196 2084 -1194
rect 2095 -1194 2102 -1190
rect 2091 -1196 2102 -1194
rect 2105 -1194 2114 -1190
rect 2105 -1196 2118 -1194
rect 2128 -1194 2137 -1190
rect 2124 -1196 2137 -1194
rect 2140 -1194 2147 -1190
rect 2140 -1196 2151 -1194
rect 2160 -1194 2169 -1190
rect 2156 -1196 2169 -1194
rect 2172 -1194 2179 -1190
rect 2172 -1196 2183 -1194
rect 2192 -1194 2200 -1190
rect 2188 -1196 2200 -1194
rect 2203 -1194 2211 -1190
rect 2203 -1196 2215 -1194
rect 2224 -1194 2233 -1190
rect 2220 -1196 2233 -1194
rect 2236 -1194 2243 -1190
rect 2236 -1196 2247 -1194
rect 2089 -1404 2093 -1399
rect 2084 -1408 2093 -1404
rect 2097 -1404 2103 -1399
rect 2097 -1408 2108 -1404
rect 2120 -1404 2125 -1399
rect 2115 -1408 2125 -1404
rect 2129 -1404 2134 -1399
rect 2129 -1408 2139 -1404
rect 2153 -1404 2159 -1399
rect 2148 -1408 2159 -1404
rect 2163 -1404 2167 -1399
rect 2163 -1408 2172 -1404
rect 2274 -1413 2286 -1409
rect 2270 -1420 2286 -1413
rect 2290 -1413 2306 -1409
rect 2290 -1420 2310 -1413
rect 2318 -1413 2332 -1409
rect 2314 -1420 2332 -1413
rect 2336 -1413 2350 -1409
rect 2336 -1420 2354 -1413
rect 2362 -1413 2377 -1409
rect 2358 -1420 2377 -1413
rect 2381 -1413 2394 -1409
rect 2381 -1420 2398 -1413
rect 2406 -1413 2420 -1409
rect 2402 -1420 2420 -1413
rect 2424 -1413 2438 -1409
rect 2424 -1420 2442 -1413
rect 2450 -1413 2465 -1409
rect 2446 -1420 2465 -1413
rect 2469 -1413 2482 -1409
rect 2469 -1420 2486 -1413
rect 2494 -1413 2508 -1409
rect 2490 -1420 2508 -1413
rect 2512 -1413 2526 -1409
rect 2512 -1420 2530 -1413
rect 2646 -1412 2658 -1408
rect 2642 -1419 2658 -1412
rect 2662 -1412 2678 -1408
rect 2662 -1419 2682 -1412
rect 2690 -1412 2704 -1408
rect 2686 -1419 2704 -1412
rect 2708 -1412 2722 -1408
rect 2708 -1419 2726 -1412
rect 2734 -1412 2749 -1408
rect 2730 -1419 2749 -1412
rect 2753 -1412 2766 -1408
rect 2753 -1419 2770 -1412
rect 2778 -1412 2792 -1408
rect 2774 -1419 2792 -1412
rect 2796 -1412 2810 -1408
rect 2796 -1419 2814 -1412
rect 2822 -1412 2837 -1408
rect 2818 -1419 2837 -1412
rect 2841 -1412 2854 -1408
rect 2841 -1419 2858 -1412
rect 2866 -1412 2880 -1408
rect 2862 -1419 2880 -1412
rect 2884 -1412 2898 -1408
rect 2884 -1419 2902 -1412
rect 3020 -1412 3032 -1408
rect 3016 -1419 3032 -1412
rect 3036 -1412 3052 -1408
rect 3036 -1419 3056 -1412
rect 3064 -1412 3078 -1408
rect 3060 -1419 3078 -1412
rect 3082 -1412 3096 -1408
rect 3082 -1419 3100 -1412
rect 3108 -1412 3123 -1408
rect 3104 -1419 3123 -1412
rect 3127 -1412 3140 -1408
rect 3127 -1419 3144 -1412
rect 3152 -1412 3166 -1408
rect 3148 -1419 3166 -1412
rect 3170 -1412 3184 -1408
rect 3170 -1419 3188 -1412
rect 3196 -1412 3211 -1408
rect 3192 -1419 3211 -1412
rect 3215 -1412 3228 -1408
rect 3215 -1419 3232 -1412
rect 3240 -1412 3254 -1408
rect 3236 -1419 3254 -1412
rect 3258 -1412 3272 -1408
rect 3258 -1419 3276 -1412
rect 3480 -1464 3488 -1460
rect 3476 -1469 3488 -1464
rect 3492 -1464 3501 -1460
rect 3492 -1469 3505 -1464
rect 3514 -1464 3523 -1460
rect 3510 -1469 3523 -1464
rect 3527 -1464 3535 -1460
rect 3527 -1469 3539 -1464
rect 3547 -1464 3556 -1460
rect 3543 -1469 3556 -1464
rect 3560 -1464 3568 -1460
rect 3560 -1469 3572 -1464
rect 3580 -1464 3589 -1460
rect 3576 -1469 3589 -1464
rect 3593 -1464 3601 -1460
rect 3593 -1469 3605 -1464
rect 3613 -1464 3622 -1460
rect 3609 -1469 3622 -1464
rect 3626 -1464 3634 -1460
rect 3626 -1469 3638 -1464
rect 2108 -1529 2128 -1525
rect 2104 -1535 2128 -1529
rect 2132 -1529 2152 -1525
rect 2132 -1535 2156 -1529
rect 2305 -1575 2325 -1571
rect 2301 -1581 2325 -1575
rect 2329 -1575 2349 -1571
rect 2329 -1581 2353 -1575
rect 2713 -1599 2733 -1595
rect 2709 -1605 2733 -1599
rect 2737 -1599 2757 -1595
rect 2737 -1605 2761 -1599
rect 3140 -1598 3160 -1594
rect 3136 -1604 3160 -1598
rect 3164 -1598 3184 -1594
rect 3164 -1604 3188 -1598
<< ndcontact >>
rect 494 1965 498 1969
rect 515 1965 519 1969
rect 523 1965 527 1969
rect 544 1965 548 1969
rect 552 1965 556 1969
rect 573 1965 577 1969
rect 581 1965 585 1969
rect 602 1965 606 1969
rect 610 1965 614 1969
rect 631 1965 635 1969
rect 639 1965 643 1969
rect 660 1965 664 1969
rect 712 1965 716 1969
rect 733 1965 737 1969
rect 741 1965 745 1969
rect 762 1965 766 1969
rect 770 1965 774 1969
rect 791 1965 795 1969
rect 799 1965 803 1969
rect 820 1965 824 1969
rect 828 1965 832 1969
rect 849 1965 853 1969
rect 857 1965 861 1969
rect 878 1965 882 1969
rect 945 1967 949 1971
rect 966 1967 970 1971
rect 974 1967 978 1971
rect 995 1967 999 1971
rect 1003 1967 1007 1971
rect 1024 1967 1028 1971
rect 1032 1967 1036 1971
rect 1053 1967 1057 1971
rect 1061 1967 1065 1971
rect 1082 1967 1086 1971
rect 1090 1967 1094 1971
rect 1111 1967 1115 1971
rect 1205 1968 1209 1972
rect 1226 1968 1230 1972
rect 1234 1968 1238 1972
rect 1255 1968 1259 1972
rect 1263 1968 1267 1972
rect 1284 1968 1288 1972
rect 1292 1968 1296 1972
rect 1313 1968 1317 1972
rect 1321 1968 1325 1972
rect 1342 1968 1346 1972
rect 1350 1968 1354 1972
rect 1371 1968 1375 1972
rect 750 1780 755 1785
rect 769 1780 774 1785
rect 781 1780 786 1785
rect 800 1780 805 1785
rect 814 1780 819 1785
rect 833 1780 838 1785
rect 926 1773 930 1777
rect 936 1773 940 1777
rect 944 1773 948 1777
rect 954 1773 958 1777
rect 963 1773 967 1777
rect 973 1773 977 1777
rect 523 1767 527 1771
rect 544 1767 548 1771
rect 552 1767 556 1771
rect 573 1767 577 1771
rect 581 1767 585 1771
rect 602 1767 606 1771
rect 610 1767 614 1771
rect 631 1767 635 1771
rect 639 1767 643 1771
rect 660 1767 664 1771
rect 668 1767 672 1771
rect 689 1767 693 1771
rect 1376 1777 1381 1782
rect 1395 1777 1400 1782
rect 1407 1777 1412 1782
rect 1426 1777 1431 1782
rect 1440 1777 1445 1782
rect 1459 1777 1464 1782
rect 1552 1770 1556 1774
rect 1562 1770 1566 1774
rect 1570 1770 1574 1774
rect 1580 1770 1584 1774
rect 1589 1770 1593 1774
rect 1599 1770 1603 1774
rect 1149 1764 1153 1768
rect 1170 1764 1174 1768
rect 1178 1764 1182 1768
rect 1199 1764 1203 1768
rect 1207 1764 1211 1768
rect 1228 1764 1232 1768
rect 1236 1764 1240 1768
rect 1257 1764 1261 1768
rect 1265 1764 1269 1768
rect 1286 1764 1290 1768
rect 1294 1764 1298 1768
rect 1315 1764 1319 1768
rect 1976 1777 1981 1782
rect 1995 1777 2000 1782
rect 2007 1777 2012 1782
rect 2026 1777 2031 1782
rect 2040 1777 2045 1782
rect 2059 1777 2064 1782
rect 2152 1770 2156 1774
rect 2162 1770 2166 1774
rect 2170 1770 2174 1774
rect 2180 1770 2184 1774
rect 2189 1770 2193 1774
rect 2199 1770 2203 1774
rect 2579 1780 2584 1785
rect 2598 1780 2603 1785
rect 2610 1780 2615 1785
rect 2629 1780 2634 1785
rect 2643 1780 2648 1785
rect 2662 1780 2667 1785
rect 2755 1773 2759 1777
rect 2765 1773 2769 1777
rect 2773 1773 2777 1777
rect 2783 1773 2787 1777
rect 2792 1773 2796 1777
rect 2802 1773 2806 1777
rect 1749 1764 1753 1768
rect 1770 1764 1774 1768
rect 1778 1764 1782 1768
rect 1799 1764 1803 1768
rect 1807 1764 1811 1768
rect 1828 1764 1832 1768
rect 1836 1764 1840 1768
rect 1857 1764 1861 1768
rect 1865 1764 1869 1768
rect 1886 1764 1890 1768
rect 1894 1764 1898 1768
rect 1915 1764 1919 1768
rect 2352 1767 2356 1771
rect 2373 1767 2377 1771
rect 2381 1767 2385 1771
rect 2402 1767 2406 1771
rect 2410 1767 2414 1771
rect 2431 1767 2435 1771
rect 2439 1767 2443 1771
rect 2460 1767 2464 1771
rect 2468 1767 2472 1771
rect 2489 1767 2493 1771
rect 2497 1767 2501 1771
rect 2518 1767 2522 1771
rect 766 1641 771 1646
rect 785 1641 790 1646
rect 797 1641 802 1646
rect 816 1641 821 1646
rect 830 1641 835 1646
rect 849 1641 854 1646
rect 1392 1638 1397 1643
rect 1411 1638 1416 1643
rect 1423 1638 1428 1643
rect 1442 1638 1447 1643
rect 1456 1638 1461 1643
rect 1475 1638 1480 1643
rect 1992 1638 1997 1643
rect 2011 1638 2016 1643
rect 2023 1638 2028 1643
rect 2042 1638 2047 1643
rect 2056 1638 2061 1643
rect 2075 1638 2080 1643
rect 2595 1641 2600 1646
rect 2614 1641 2619 1646
rect 2626 1641 2631 1646
rect 2645 1641 2650 1646
rect 2659 1641 2664 1646
rect 2678 1641 2683 1646
rect 533 1511 537 1515
rect 554 1511 558 1515
rect 562 1511 566 1515
rect 583 1511 587 1515
rect 591 1511 595 1515
rect 612 1511 616 1515
rect 620 1511 624 1515
rect 641 1511 645 1515
rect 649 1511 653 1515
rect 670 1511 674 1515
rect 678 1511 682 1515
rect 699 1511 703 1515
rect 1159 1508 1163 1512
rect 1180 1508 1184 1512
rect 1188 1508 1192 1512
rect 1209 1508 1213 1512
rect 1217 1508 1221 1512
rect 1238 1508 1242 1512
rect 1246 1508 1250 1512
rect 1267 1508 1271 1512
rect 1275 1508 1279 1512
rect 1296 1508 1300 1512
rect 1304 1508 1308 1512
rect 1325 1508 1329 1512
rect 1759 1508 1763 1512
rect 1780 1508 1784 1512
rect 1788 1508 1792 1512
rect 1809 1508 1813 1512
rect 1817 1508 1821 1512
rect 1838 1508 1842 1512
rect 1846 1508 1850 1512
rect 1867 1508 1871 1512
rect 1875 1508 1879 1512
rect 1896 1508 1900 1512
rect 1904 1508 1908 1512
rect 1925 1508 1929 1512
rect 2362 1511 2366 1515
rect 2383 1511 2387 1515
rect 2391 1511 2395 1515
rect 2412 1511 2416 1515
rect 2420 1511 2424 1515
rect 2441 1511 2445 1515
rect 2449 1511 2453 1515
rect 2470 1511 2474 1515
rect 2478 1511 2482 1515
rect 2499 1511 2503 1515
rect 2507 1511 2511 1515
rect 2528 1511 2532 1515
rect 547 1150 551 1154
rect 568 1150 572 1154
rect 576 1150 580 1154
rect 597 1150 601 1154
rect 605 1150 609 1154
rect 626 1150 630 1154
rect 634 1150 638 1154
rect 655 1150 659 1154
rect 663 1150 667 1154
rect 684 1150 688 1154
rect 692 1150 696 1154
rect 713 1150 717 1154
rect 765 1150 769 1154
rect 786 1150 790 1154
rect 794 1150 798 1154
rect 815 1150 819 1154
rect 823 1150 827 1154
rect 844 1150 848 1154
rect 852 1150 856 1154
rect 873 1150 877 1154
rect 881 1150 885 1154
rect 902 1150 906 1154
rect 910 1150 914 1154
rect 931 1150 935 1154
rect 998 1152 1002 1156
rect 1019 1152 1023 1156
rect 1027 1152 1031 1156
rect 1048 1152 1052 1156
rect 1056 1152 1060 1156
rect 1077 1152 1081 1156
rect 1085 1152 1089 1156
rect 1106 1152 1110 1156
rect 1114 1152 1118 1156
rect 1135 1152 1139 1156
rect 1143 1152 1147 1156
rect 1164 1152 1168 1156
rect 1258 1153 1262 1157
rect 1279 1153 1283 1157
rect 1287 1153 1291 1157
rect 1308 1153 1312 1157
rect 1316 1153 1320 1157
rect 1337 1153 1341 1157
rect 1345 1153 1349 1157
rect 1366 1153 1370 1157
rect 1374 1153 1378 1157
rect 1395 1153 1399 1157
rect 1403 1153 1407 1157
rect 1424 1153 1428 1157
rect -410 1013 -405 1018
rect -391 1013 -386 1018
rect -379 1013 -374 1018
rect -360 1013 -355 1018
rect -346 1013 -341 1018
rect -327 1013 -322 1018
rect -274 1014 -269 1019
rect -255 1014 -250 1019
rect -243 1014 -238 1019
rect -224 1014 -219 1019
rect -210 1014 -205 1019
rect -191 1014 -186 1019
rect -139 1015 -134 1020
rect -120 1015 -115 1020
rect -108 1015 -103 1020
rect -89 1015 -84 1020
rect -75 1015 -70 1020
rect -56 1015 -51 1020
rect -2 1013 3 1018
rect 17 1013 22 1018
rect 29 1013 34 1018
rect 48 1013 53 1018
rect 62 1013 67 1018
rect 81 1013 86 1018
rect 803 965 808 970
rect 822 965 827 970
rect 834 965 839 970
rect 853 965 858 970
rect 867 965 872 970
rect 886 965 891 970
rect 979 958 983 962
rect 989 958 993 962
rect 997 958 1001 962
rect 1007 958 1011 962
rect 1016 958 1020 962
rect 1026 958 1030 962
rect 576 952 580 956
rect -411 893 -406 898
rect -392 893 -387 898
rect -380 893 -375 898
rect -361 893 -356 898
rect -347 893 -342 898
rect -328 893 -323 898
rect -265 894 -260 899
rect -246 894 -241 899
rect -234 894 -229 899
rect -215 894 -210 899
rect -201 894 -196 899
rect -182 894 -177 899
rect -135 897 -130 902
rect -116 897 -111 902
rect -104 897 -99 902
rect -85 897 -80 902
rect -71 897 -66 902
rect -52 897 -47 902
rect 597 952 601 956
rect 605 952 609 956
rect 626 952 630 956
rect 634 952 638 956
rect 655 952 659 956
rect 663 952 667 956
rect 684 952 688 956
rect 692 952 696 956
rect 713 952 717 956
rect 721 952 725 956
rect 742 952 746 956
rect 1429 962 1434 967
rect 1448 962 1453 967
rect 1460 962 1465 967
rect 1479 962 1484 967
rect 1493 962 1498 967
rect 1512 962 1517 967
rect 1605 955 1609 959
rect 1615 955 1619 959
rect 1623 955 1627 959
rect 1633 955 1637 959
rect 1642 955 1646 959
rect 1652 955 1656 959
rect 1202 949 1206 953
rect 1223 949 1227 953
rect 1231 949 1235 953
rect 1252 949 1256 953
rect 1260 949 1264 953
rect 1281 949 1285 953
rect 1289 949 1293 953
rect 1310 949 1314 953
rect 1318 949 1322 953
rect 1339 949 1343 953
rect 1347 949 1351 953
rect 1368 949 1372 953
rect 2029 962 2034 967
rect 2048 962 2053 967
rect 2060 962 2065 967
rect 2079 962 2084 967
rect 2093 962 2098 967
rect 2112 962 2117 967
rect 2205 955 2209 959
rect 2215 955 2219 959
rect 2223 955 2227 959
rect 2233 955 2237 959
rect 2242 955 2246 959
rect 2252 955 2256 959
rect 2632 965 2637 970
rect 2651 965 2656 970
rect 2663 965 2668 970
rect 2682 965 2687 970
rect 2696 965 2701 970
rect 2715 965 2720 970
rect 2808 958 2812 962
rect 2818 958 2822 962
rect 2826 958 2830 962
rect 2836 958 2840 962
rect 2845 958 2849 962
rect 2855 958 2859 962
rect 1802 949 1806 953
rect 1823 949 1827 953
rect 1831 949 1835 953
rect 1852 949 1856 953
rect 1860 949 1864 953
rect 1881 949 1885 953
rect 1889 949 1893 953
rect 1910 949 1914 953
rect 1918 949 1922 953
rect 1939 949 1943 953
rect 1947 949 1951 953
rect 1968 949 1972 953
rect 2405 952 2409 956
rect 2426 952 2430 956
rect 2434 952 2438 956
rect 2455 952 2459 956
rect 2463 952 2467 956
rect 2484 952 2488 956
rect 2492 952 2496 956
rect 2513 952 2517 956
rect 2521 952 2525 956
rect 2542 952 2546 956
rect 2550 952 2554 956
rect 2571 952 2575 956
rect 6 896 11 901
rect 25 896 30 901
rect 37 896 42 901
rect 56 896 61 901
rect 70 896 75 901
rect 89 896 94 901
rect 819 826 824 831
rect 838 826 843 831
rect 850 826 855 831
rect 869 826 874 831
rect 883 826 888 831
rect 902 826 907 831
rect 1445 823 1450 828
rect 1464 823 1469 828
rect 1476 823 1481 828
rect 1495 823 1500 828
rect 1509 823 1514 828
rect 1528 823 1533 828
rect 2045 823 2050 828
rect 2064 823 2069 828
rect 2076 823 2081 828
rect 2095 823 2100 828
rect 2109 823 2114 828
rect 2128 823 2133 828
rect 2648 826 2653 831
rect 2667 826 2672 831
rect 2679 826 2684 831
rect 2698 826 2703 831
rect 2712 826 2717 831
rect 2731 826 2736 831
rect 586 696 590 700
rect 607 696 611 700
rect 615 696 619 700
rect 636 696 640 700
rect 644 696 648 700
rect 665 696 669 700
rect 673 696 677 700
rect 694 696 698 700
rect 702 696 706 700
rect 723 696 727 700
rect 731 696 735 700
rect 752 696 756 700
rect 1212 693 1216 697
rect 1233 693 1237 697
rect 1241 693 1245 697
rect 1262 693 1266 697
rect 1270 693 1274 697
rect 1291 693 1295 697
rect 1299 693 1303 697
rect 1320 693 1324 697
rect 1328 693 1332 697
rect 1349 693 1353 697
rect 1357 693 1361 697
rect 1378 693 1382 697
rect 1812 693 1816 697
rect 1833 693 1837 697
rect 1841 693 1845 697
rect 1862 693 1866 697
rect 1870 693 1874 697
rect 1891 693 1895 697
rect 1899 693 1903 697
rect 1920 693 1924 697
rect 1928 693 1932 697
rect 1949 693 1953 697
rect 1957 693 1961 697
rect 1978 693 1982 697
rect 2415 696 2419 700
rect 2436 696 2440 700
rect 2444 696 2448 700
rect 2465 696 2469 700
rect 2473 696 2477 700
rect 2494 696 2498 700
rect 2502 696 2506 700
rect 2523 696 2527 700
rect 2531 696 2535 700
rect 2552 696 2556 700
rect 2560 696 2564 700
rect 2581 696 2585 700
rect -391 570 -386 575
rect -372 570 -367 575
rect -360 570 -355 575
rect -341 570 -336 575
rect -327 570 -322 575
rect -308 570 -303 575
rect -255 571 -250 576
rect -236 571 -231 576
rect -224 571 -219 576
rect -205 571 -200 576
rect -191 571 -186 576
rect -172 571 -167 576
rect -120 572 -115 577
rect -101 572 -96 577
rect -89 572 -84 577
rect -70 572 -65 577
rect -56 572 -51 577
rect -37 572 -32 577
rect 17 570 22 575
rect 36 570 41 575
rect 48 570 53 575
rect 67 570 72 575
rect 81 570 86 575
rect 100 570 105 575
rect -392 450 -387 455
rect -373 450 -368 455
rect -361 450 -356 455
rect -342 450 -337 455
rect -328 450 -323 455
rect -309 450 -304 455
rect -246 451 -241 456
rect -227 451 -222 456
rect -215 451 -210 456
rect -196 451 -191 456
rect -182 451 -177 456
rect -163 451 -158 456
rect -116 454 -111 459
rect -97 454 -92 459
rect -85 454 -80 459
rect -66 454 -61 459
rect -52 454 -47 459
rect -33 454 -28 459
rect 25 453 30 458
rect 44 453 49 458
rect 56 453 61 458
rect 75 453 80 458
rect 89 453 94 458
rect 108 453 113 458
rect -1052 396 -1047 401
rect -1033 396 -1028 401
rect -1021 396 -1016 401
rect -1002 396 -997 401
rect -988 396 -983 401
rect -969 396 -964 401
rect -1239 388 -1235 392
rect -1191 388 -1187 392
rect -1050 295 -1045 300
rect -1031 295 -1026 300
rect -1019 295 -1014 300
rect -1000 295 -995 300
rect -986 295 -981 300
rect -967 295 -962 300
rect -1047 196 -1042 201
rect -1028 196 -1023 201
rect -1016 196 -1011 201
rect -997 196 -992 201
rect -983 196 -978 201
rect -964 196 -959 201
rect -1241 169 -1237 173
rect -1193 169 -1189 173
rect -378 145 -373 150
rect -359 145 -354 150
rect -347 145 -342 150
rect -328 145 -323 150
rect -314 145 -309 150
rect -295 145 -290 150
rect -242 146 -237 151
rect -223 146 -218 151
rect -211 146 -206 151
rect -192 146 -187 151
rect -178 146 -173 151
rect -159 146 -154 151
rect -107 147 -102 152
rect -88 147 -83 152
rect -76 147 -71 152
rect -57 147 -52 152
rect -43 147 -38 152
rect -24 147 -19 152
rect 30 145 35 150
rect 49 145 54 150
rect 61 145 66 150
rect 80 145 85 150
rect 94 145 99 150
rect 113 145 118 150
rect -1045 88 -1040 93
rect -1026 88 -1021 93
rect -1014 88 -1009 93
rect -995 88 -990 93
rect -981 88 -976 93
rect -962 88 -957 93
rect -379 25 -374 30
rect -360 25 -355 30
rect -348 25 -343 30
rect -329 25 -324 30
rect -315 25 -310 30
rect -296 25 -291 30
rect -233 26 -228 31
rect -214 26 -209 31
rect -202 26 -197 31
rect -183 26 -178 31
rect -169 26 -164 31
rect -150 26 -145 31
rect -103 29 -98 34
rect -84 29 -79 34
rect -72 29 -67 34
rect -53 29 -48 34
rect -39 29 -34 34
rect -20 29 -15 34
rect 38 28 43 33
rect 57 28 62 33
rect 69 28 74 33
rect 88 28 93 33
rect 102 28 107 33
rect 121 28 126 33
rect 2077 -28 2081 -24
rect 2125 -28 2129 -24
rect 2602 -27 2606 -23
rect 2347 -33 2351 -29
rect 2395 -33 2399 -29
rect 2650 -27 2654 -23
rect 2870 -27 2874 -23
rect 2918 -27 2922 -23
rect -326 -305 -321 -300
rect -307 -305 -302 -300
rect -295 -305 -290 -300
rect -276 -305 -271 -300
rect -262 -305 -257 -300
rect -243 -305 -238 -300
rect -190 -304 -185 -299
rect -171 -304 -166 -299
rect -159 -304 -154 -299
rect -140 -304 -135 -299
rect -126 -304 -121 -299
rect -107 -304 -102 -299
rect -55 -303 -50 -298
rect -36 -303 -31 -298
rect -24 -303 -19 -298
rect -5 -303 0 -298
rect 9 -303 14 -298
rect 28 -303 33 -298
rect 82 -305 87 -300
rect 101 -305 106 -300
rect 113 -305 118 -300
rect 132 -305 137 -300
rect 146 -305 151 -300
rect 165 -305 170 -300
rect 3426 -219 3430 -215
rect 3451 -219 3455 -215
rect 3460 -219 3464 -215
rect 3485 -219 3489 -215
rect 3493 -219 3497 -215
rect 3518 -219 3522 -215
rect 3526 -219 3530 -215
rect 3551 -219 3555 -215
rect 3559 -219 3563 -215
rect 3584 -219 3588 -215
rect 2219 -290 2223 -286
rect 2255 -290 2259 -286
rect 2263 -290 2267 -286
rect 2299 -290 2303 -286
rect 2307 -290 2311 -286
rect 2343 -290 2347 -286
rect 2351 -290 2355 -286
rect 2387 -290 2391 -286
rect 2395 -290 2399 -286
rect 2431 -290 2435 -286
rect 2439 -290 2443 -286
rect 2475 -290 2479 -286
rect 2601 -290 2605 -286
rect 2637 -290 2641 -286
rect 2645 -290 2649 -286
rect 2681 -290 2685 -286
rect 2689 -290 2693 -286
rect 2725 -290 2729 -286
rect 2733 -290 2737 -286
rect 2769 -290 2773 -286
rect 2777 -290 2781 -286
rect 2813 -290 2817 -286
rect 2821 -290 2825 -286
rect 2857 -290 2861 -286
rect 2983 -290 2987 -286
rect 3019 -290 3023 -286
rect 3027 -290 3031 -286
rect 3063 -290 3067 -286
rect 3071 -290 3075 -286
rect 3107 -290 3111 -286
rect 3115 -290 3119 -286
rect 3151 -290 3155 -286
rect 3159 -290 3163 -286
rect 3195 -290 3199 -286
rect 3203 -290 3207 -286
rect 3239 -290 3243 -286
rect 2041 -317 2046 -312
rect 2060 -317 2065 -312
rect 2072 -317 2077 -312
rect 2091 -317 2096 -312
rect 2105 -317 2110 -312
rect 2124 -317 2129 -312
rect -327 -425 -322 -420
rect -308 -425 -303 -420
rect -296 -425 -291 -420
rect -277 -425 -272 -420
rect -263 -425 -258 -420
rect -244 -425 -239 -420
rect -181 -424 -176 -419
rect -162 -424 -157 -419
rect -150 -424 -145 -419
rect -131 -424 -126 -419
rect -117 -424 -112 -419
rect -98 -424 -93 -419
rect -51 -421 -46 -416
rect -32 -421 -27 -416
rect -20 -421 -15 -416
rect -1 -421 4 -416
rect 13 -421 18 -416
rect 32 -421 37 -416
rect 90 -422 95 -417
rect 109 -422 114 -417
rect 121 -422 126 -417
rect 140 -422 145 -417
rect 154 -422 159 -417
rect 173 -422 178 -417
rect 401 -485 406 -480
rect 420 -485 425 -480
rect 432 -485 437 -480
rect 451 -485 456 -480
rect 465 -485 470 -480
rect 484 -485 489 -480
rect -270 -591 -265 -586
rect -251 -591 -246 -586
rect -239 -591 -234 -586
rect -220 -591 -215 -586
rect -206 -591 -201 -586
rect -187 -591 -182 -586
rect 2057 -603 2061 -599
rect -94 -647 -89 -642
rect -75 -647 -70 -642
rect -63 -647 -58 -642
rect -44 -647 -39 -642
rect -30 -647 -25 -642
rect -11 -647 -6 -642
rect 2080 -603 2084 -599
rect 2091 -603 2095 -599
rect 2114 -603 2118 -599
rect 2124 -603 2128 -599
rect 2147 -603 2151 -599
rect 2156 -603 2160 -599
rect 2179 -603 2183 -599
rect 2188 -603 2192 -599
rect 2211 -603 2215 -599
rect 2220 -603 2224 -599
rect 2243 -603 2247 -599
rect 160 -657 165 -652
rect 179 -657 184 -652
rect 191 -657 196 -652
rect 210 -657 215 -652
rect 224 -657 229 -652
rect 243 -657 248 -652
rect 2056 -850 2060 -846
rect 2079 -850 2083 -846
rect 2090 -850 2094 -846
rect 2113 -850 2117 -846
rect 2123 -850 2127 -846
rect 2146 -850 2150 -846
rect 2155 -850 2159 -846
rect 2178 -850 2182 -846
rect 2187 -850 2191 -846
rect 2210 -850 2214 -846
rect 2219 -850 2223 -846
rect 2242 -850 2246 -846
rect 2410 -910 2414 -906
rect 2446 -910 2450 -906
rect 2454 -910 2458 -906
rect 2490 -910 2494 -906
rect 2498 -910 2502 -906
rect 2534 -910 2538 -906
rect 2542 -910 2546 -906
rect 2578 -910 2582 -906
rect 2586 -910 2590 -906
rect 2622 -910 2626 -906
rect 2630 -910 2634 -906
rect 2666 -910 2670 -906
rect 2060 -1076 2064 -1072
rect 2083 -1076 2087 -1072
rect 2094 -1076 2098 -1072
rect 2117 -1076 2121 -1072
rect 2127 -1076 2131 -1072
rect 2150 -1076 2154 -1072
rect 2159 -1076 2163 -1072
rect 2182 -1076 2186 -1072
rect 2191 -1076 2195 -1072
rect 2214 -1076 2218 -1072
rect 2223 -1076 2227 -1072
rect 2246 -1076 2250 -1072
rect 2057 -1283 2061 -1279
rect 2080 -1283 2084 -1279
rect 2091 -1283 2095 -1279
rect 2114 -1283 2118 -1279
rect 2124 -1283 2128 -1279
rect 2147 -1283 2151 -1279
rect 2156 -1283 2160 -1279
rect 2179 -1283 2183 -1279
rect 2188 -1283 2192 -1279
rect 2211 -1283 2215 -1279
rect 2220 -1283 2224 -1279
rect 2243 -1283 2247 -1279
rect 2084 -1462 2089 -1457
rect 2103 -1462 2108 -1457
rect 2115 -1462 2120 -1457
rect 2134 -1462 2139 -1457
rect 2148 -1462 2153 -1457
rect 2167 -1462 2172 -1457
rect 2270 -1516 2274 -1512
rect 2306 -1516 2310 -1512
rect 2314 -1516 2318 -1512
rect 2350 -1516 2354 -1512
rect 2358 -1516 2362 -1512
rect 2394 -1516 2398 -1512
rect 2402 -1516 2406 -1512
rect 2438 -1516 2442 -1512
rect 2446 -1516 2450 -1512
rect 2482 -1516 2486 -1512
rect 2490 -1516 2494 -1512
rect 2526 -1516 2530 -1512
rect 2642 -1515 2646 -1511
rect 2678 -1515 2682 -1511
rect 2686 -1515 2690 -1511
rect 2722 -1515 2726 -1511
rect 2730 -1515 2734 -1511
rect 2766 -1515 2770 -1511
rect 2774 -1515 2778 -1511
rect 2810 -1515 2814 -1511
rect 2818 -1515 2822 -1511
rect 2854 -1515 2858 -1511
rect 2862 -1515 2866 -1511
rect 2898 -1515 2902 -1511
rect 3016 -1515 3020 -1511
rect 3052 -1515 3056 -1511
rect 3060 -1515 3064 -1511
rect 3096 -1515 3100 -1511
rect 3104 -1515 3108 -1511
rect 3140 -1515 3144 -1511
rect 3148 -1515 3152 -1511
rect 3184 -1515 3188 -1511
rect 3192 -1515 3196 -1511
rect 3228 -1515 3232 -1511
rect 3236 -1515 3240 -1511
rect 3272 -1515 3276 -1511
rect 3476 -1546 3480 -1542
rect 3501 -1546 3505 -1542
rect 3510 -1546 3514 -1542
rect 3535 -1546 3539 -1542
rect 3543 -1546 3547 -1542
rect 3568 -1546 3572 -1542
rect 3576 -1546 3580 -1542
rect 3601 -1546 3605 -1542
rect 3609 -1546 3613 -1542
rect 3634 -1546 3638 -1542
rect 2104 -1567 2108 -1563
rect 2152 -1567 2156 -1563
rect 2301 -1613 2305 -1609
rect 2349 -1613 2353 -1609
rect 2709 -1637 2713 -1633
rect 2757 -1637 2761 -1633
rect 3136 -1636 3140 -1632
rect 3184 -1636 3188 -1632
<< pdcontact >>
rect 494 2037 498 2041
rect 515 2037 519 2041
rect 523 2037 527 2041
rect 544 2037 548 2041
rect 552 2037 556 2041
rect 573 2037 577 2041
rect 581 2037 585 2041
rect 602 2037 606 2041
rect 610 2037 614 2041
rect 631 2037 635 2041
rect 639 2037 643 2041
rect 660 2037 664 2041
rect 712 2037 716 2041
rect 733 2037 737 2041
rect 741 2037 745 2041
rect 762 2037 766 2041
rect 770 2037 774 2041
rect 791 2037 795 2041
rect 799 2037 803 2041
rect 820 2037 824 2041
rect 828 2037 832 2041
rect 849 2037 853 2041
rect 857 2037 861 2041
rect 878 2037 882 2041
rect 945 2039 949 2043
rect 966 2039 970 2043
rect 974 2039 978 2043
rect 995 2039 999 2043
rect 1003 2039 1007 2043
rect 1024 2039 1028 2043
rect 1032 2039 1036 2043
rect 1053 2039 1057 2043
rect 1061 2039 1065 2043
rect 1082 2039 1086 2043
rect 1090 2039 1094 2043
rect 1111 2039 1115 2043
rect 1205 2040 1209 2044
rect 1226 2040 1230 2044
rect 1234 2040 1238 2044
rect 1255 2040 1259 2044
rect 1263 2040 1267 2044
rect 1284 2040 1288 2044
rect 1292 2040 1296 2044
rect 1313 2040 1317 2044
rect 1321 2040 1325 2044
rect 1342 2040 1346 2044
rect 1350 2040 1354 2044
rect 1371 2040 1375 2044
rect 523 1839 527 1843
rect 544 1839 548 1843
rect 552 1839 556 1843
rect 573 1839 577 1843
rect 581 1839 585 1843
rect 602 1839 606 1843
rect 610 1839 614 1843
rect 631 1839 635 1843
rect 639 1839 643 1843
rect 660 1839 664 1843
rect 668 1839 672 1843
rect 689 1839 693 1843
rect 750 1838 755 1843
rect 769 1838 774 1843
rect 781 1838 786 1843
rect 800 1838 805 1843
rect 814 1838 819 1843
rect 833 1838 838 1843
rect 1149 1836 1153 1840
rect 1170 1836 1174 1840
rect 1178 1836 1182 1840
rect 1199 1836 1203 1840
rect 1207 1836 1211 1840
rect 1228 1836 1232 1840
rect 1236 1836 1240 1840
rect 1257 1836 1261 1840
rect 1265 1836 1269 1840
rect 1286 1836 1290 1840
rect 1294 1836 1298 1840
rect 1315 1836 1319 1840
rect 1376 1835 1381 1840
rect 926 1814 930 1818
rect 936 1814 940 1818
rect 944 1814 948 1818
rect 954 1814 958 1818
rect 963 1814 967 1818
rect 973 1814 977 1818
rect 1395 1835 1400 1840
rect 1407 1835 1412 1840
rect 1426 1835 1431 1840
rect 1440 1835 1445 1840
rect 1459 1835 1464 1840
rect 1749 1836 1753 1840
rect 1770 1836 1774 1840
rect 1778 1836 1782 1840
rect 1799 1836 1803 1840
rect 1807 1836 1811 1840
rect 1828 1836 1832 1840
rect 1836 1836 1840 1840
rect 1857 1836 1861 1840
rect 1865 1836 1869 1840
rect 1886 1836 1890 1840
rect 1894 1836 1898 1840
rect 1915 1836 1919 1840
rect 1976 1835 1981 1840
rect 1552 1811 1556 1815
rect 1562 1811 1566 1815
rect 1570 1811 1574 1815
rect 1580 1811 1584 1815
rect 1589 1811 1593 1815
rect 1599 1811 1603 1815
rect 1995 1835 2000 1840
rect 2007 1835 2012 1840
rect 2026 1835 2031 1840
rect 2040 1835 2045 1840
rect 2059 1835 2064 1840
rect 2352 1839 2356 1843
rect 2373 1839 2377 1843
rect 2381 1839 2385 1843
rect 2402 1839 2406 1843
rect 2410 1839 2414 1843
rect 2431 1839 2435 1843
rect 2439 1839 2443 1843
rect 2460 1839 2464 1843
rect 2468 1839 2472 1843
rect 2489 1839 2493 1843
rect 2497 1839 2501 1843
rect 2518 1839 2522 1843
rect 2579 1838 2584 1843
rect 2152 1811 2156 1815
rect 2162 1811 2166 1815
rect 2170 1811 2174 1815
rect 2180 1811 2184 1815
rect 2189 1811 2193 1815
rect 2199 1811 2203 1815
rect 2598 1838 2603 1843
rect 2610 1838 2615 1843
rect 2629 1838 2634 1843
rect 2643 1838 2648 1843
rect 2662 1838 2667 1843
rect 2755 1814 2759 1818
rect 2765 1814 2769 1818
rect 2773 1814 2777 1818
rect 2783 1814 2787 1818
rect 2792 1814 2796 1818
rect 2802 1814 2806 1818
rect 766 1699 771 1704
rect 785 1699 790 1704
rect 797 1699 802 1704
rect 816 1699 821 1704
rect 830 1699 835 1704
rect 849 1699 854 1704
rect 1392 1696 1397 1701
rect 1411 1696 1416 1701
rect 1423 1696 1428 1701
rect 1442 1696 1447 1701
rect 1456 1696 1461 1701
rect 1475 1696 1480 1701
rect 1992 1696 1997 1701
rect 2011 1696 2016 1701
rect 2023 1696 2028 1701
rect 2042 1696 2047 1701
rect 2056 1696 2061 1701
rect 2075 1696 2080 1701
rect 2595 1699 2600 1704
rect 2614 1699 2619 1704
rect 2626 1699 2631 1704
rect 2645 1699 2650 1704
rect 2659 1699 2664 1704
rect 2678 1699 2683 1704
rect 533 1583 537 1587
rect 554 1583 558 1587
rect 562 1583 566 1587
rect 583 1583 587 1587
rect 591 1583 595 1587
rect 612 1583 616 1587
rect 620 1583 624 1587
rect 641 1583 645 1587
rect 649 1583 653 1587
rect 670 1583 674 1587
rect 678 1583 682 1587
rect 699 1583 703 1587
rect 1159 1580 1163 1584
rect 1180 1580 1184 1584
rect 1188 1580 1192 1584
rect 1209 1580 1213 1584
rect 1217 1580 1221 1584
rect 1238 1580 1242 1584
rect 1246 1580 1250 1584
rect 1267 1580 1271 1584
rect 1275 1580 1279 1584
rect 1296 1580 1300 1584
rect 1304 1580 1308 1584
rect 1325 1580 1329 1584
rect 1759 1580 1763 1584
rect 1780 1580 1784 1584
rect 1788 1580 1792 1584
rect 1809 1580 1813 1584
rect 1817 1580 1821 1584
rect 1838 1580 1842 1584
rect 1846 1580 1850 1584
rect 1867 1580 1871 1584
rect 1875 1580 1879 1584
rect 1896 1580 1900 1584
rect 1904 1580 1908 1584
rect 1925 1580 1929 1584
rect 2362 1583 2366 1587
rect 2383 1583 2387 1587
rect 2391 1583 2395 1587
rect 2412 1583 2416 1587
rect 2420 1583 2424 1587
rect 2441 1583 2445 1587
rect 2449 1583 2453 1587
rect 2470 1583 2474 1587
rect 2478 1583 2482 1587
rect 2499 1583 2503 1587
rect 2507 1583 2511 1587
rect 2528 1583 2532 1587
rect 547 1222 551 1226
rect 568 1222 572 1226
rect 576 1222 580 1226
rect 597 1222 601 1226
rect 605 1222 609 1226
rect 626 1222 630 1226
rect 634 1222 638 1226
rect 655 1222 659 1226
rect 663 1222 667 1226
rect 684 1222 688 1226
rect 692 1222 696 1226
rect 713 1222 717 1226
rect 765 1222 769 1226
rect 786 1222 790 1226
rect 794 1222 798 1226
rect 815 1222 819 1226
rect 823 1222 827 1226
rect 844 1222 848 1226
rect 852 1222 856 1226
rect 873 1222 877 1226
rect 881 1222 885 1226
rect 902 1222 906 1226
rect 910 1222 914 1226
rect 931 1222 935 1226
rect 998 1224 1002 1228
rect 1019 1224 1023 1228
rect 1027 1224 1031 1228
rect 1048 1224 1052 1228
rect 1056 1224 1060 1228
rect 1077 1224 1081 1228
rect 1085 1224 1089 1228
rect 1106 1224 1110 1228
rect 1114 1224 1118 1228
rect 1135 1224 1139 1228
rect 1143 1224 1147 1228
rect 1164 1224 1168 1228
rect 1258 1225 1262 1229
rect 1279 1225 1283 1229
rect 1287 1225 1291 1229
rect 1308 1225 1312 1229
rect 1316 1225 1320 1229
rect 1337 1225 1341 1229
rect 1345 1225 1349 1229
rect 1366 1225 1370 1229
rect 1374 1225 1378 1229
rect 1395 1225 1399 1229
rect 1403 1225 1407 1229
rect 1424 1225 1428 1229
rect -410 1071 -405 1076
rect -391 1071 -386 1076
rect -379 1071 -374 1076
rect -360 1071 -355 1076
rect -346 1071 -341 1076
rect -327 1071 -322 1076
rect -274 1072 -269 1077
rect -255 1072 -250 1077
rect -243 1072 -238 1077
rect -224 1072 -219 1077
rect -210 1072 -205 1077
rect -191 1072 -186 1077
rect -139 1073 -134 1078
rect -120 1073 -115 1078
rect -108 1073 -103 1078
rect -89 1073 -84 1078
rect -75 1073 -70 1078
rect -56 1073 -51 1078
rect -2 1071 3 1076
rect 17 1071 22 1076
rect 29 1071 34 1076
rect 48 1071 53 1076
rect 62 1071 67 1076
rect 81 1071 86 1076
rect 576 1024 580 1028
rect 597 1024 601 1028
rect 605 1024 609 1028
rect 626 1024 630 1028
rect 634 1024 638 1028
rect 655 1024 659 1028
rect 663 1024 667 1028
rect 684 1024 688 1028
rect 692 1024 696 1028
rect 713 1024 717 1028
rect 721 1024 725 1028
rect 742 1024 746 1028
rect 803 1023 808 1028
rect -411 951 -406 956
rect -392 951 -387 956
rect -380 951 -375 956
rect -361 951 -356 956
rect -347 951 -342 956
rect -328 951 -323 956
rect -265 952 -260 957
rect -246 952 -241 957
rect -234 952 -229 957
rect -215 952 -210 957
rect -201 952 -196 957
rect -182 952 -177 957
rect -135 955 -130 960
rect -116 955 -111 960
rect -104 955 -99 960
rect -85 955 -80 960
rect -71 955 -66 960
rect -52 955 -47 960
rect 6 954 11 959
rect 25 954 30 959
rect 37 954 42 959
rect 56 954 61 959
rect 70 954 75 959
rect 89 954 94 959
rect 822 1023 827 1028
rect 834 1023 839 1028
rect 853 1023 858 1028
rect 867 1023 872 1028
rect 886 1023 891 1028
rect 1202 1021 1206 1025
rect 1223 1021 1227 1025
rect 1231 1021 1235 1025
rect 1252 1021 1256 1025
rect 1260 1021 1264 1025
rect 1281 1021 1285 1025
rect 1289 1021 1293 1025
rect 1310 1021 1314 1025
rect 1318 1021 1322 1025
rect 1339 1021 1343 1025
rect 1347 1021 1351 1025
rect 1368 1021 1372 1025
rect 1429 1020 1434 1025
rect 979 999 983 1003
rect 989 999 993 1003
rect 997 999 1001 1003
rect 1007 999 1011 1003
rect 1016 999 1020 1003
rect 1026 999 1030 1003
rect 1448 1020 1453 1025
rect 1460 1020 1465 1025
rect 1479 1020 1484 1025
rect 1493 1020 1498 1025
rect 1512 1020 1517 1025
rect 1802 1021 1806 1025
rect 1823 1021 1827 1025
rect 1831 1021 1835 1025
rect 1852 1021 1856 1025
rect 1860 1021 1864 1025
rect 1881 1021 1885 1025
rect 1889 1021 1893 1025
rect 1910 1021 1914 1025
rect 1918 1021 1922 1025
rect 1939 1021 1943 1025
rect 1947 1021 1951 1025
rect 1968 1021 1972 1025
rect 2029 1020 2034 1025
rect 1605 996 1609 1000
rect 1615 996 1619 1000
rect 1623 996 1627 1000
rect 1633 996 1637 1000
rect 1642 996 1646 1000
rect 1652 996 1656 1000
rect 2048 1020 2053 1025
rect 2060 1020 2065 1025
rect 2079 1020 2084 1025
rect 2093 1020 2098 1025
rect 2112 1020 2117 1025
rect 2405 1024 2409 1028
rect 2426 1024 2430 1028
rect 2434 1024 2438 1028
rect 2455 1024 2459 1028
rect 2463 1024 2467 1028
rect 2484 1024 2488 1028
rect 2492 1024 2496 1028
rect 2513 1024 2517 1028
rect 2521 1024 2525 1028
rect 2542 1024 2546 1028
rect 2550 1024 2554 1028
rect 2571 1024 2575 1028
rect 2632 1023 2637 1028
rect 2205 996 2209 1000
rect 2215 996 2219 1000
rect 2223 996 2227 1000
rect 2233 996 2237 1000
rect 2242 996 2246 1000
rect 2252 996 2256 1000
rect 2651 1023 2656 1028
rect 2663 1023 2668 1028
rect 2682 1023 2687 1028
rect 2696 1023 2701 1028
rect 2715 1023 2720 1028
rect 2808 999 2812 1003
rect 2818 999 2822 1003
rect 2826 999 2830 1003
rect 2836 999 2840 1003
rect 2845 999 2849 1003
rect 2855 999 2859 1003
rect 819 884 824 889
rect 838 884 843 889
rect 850 884 855 889
rect 869 884 874 889
rect 883 884 888 889
rect 902 884 907 889
rect 1445 881 1450 886
rect 1464 881 1469 886
rect 1476 881 1481 886
rect 1495 881 1500 886
rect 1509 881 1514 886
rect 1528 881 1533 886
rect 2045 881 2050 886
rect 2064 881 2069 886
rect 2076 881 2081 886
rect 2095 881 2100 886
rect 2109 881 2114 886
rect 2128 881 2133 886
rect 2648 884 2653 889
rect 2667 884 2672 889
rect 2679 884 2684 889
rect 2698 884 2703 889
rect 2712 884 2717 889
rect 2731 884 2736 889
rect 586 768 590 772
rect 607 768 611 772
rect 615 768 619 772
rect 636 768 640 772
rect 644 768 648 772
rect 665 768 669 772
rect 673 768 677 772
rect 694 768 698 772
rect 702 768 706 772
rect 723 768 727 772
rect 731 768 735 772
rect 752 768 756 772
rect 1212 765 1216 769
rect 1233 765 1237 769
rect 1241 765 1245 769
rect 1262 765 1266 769
rect 1270 765 1274 769
rect 1291 765 1295 769
rect 1299 765 1303 769
rect 1320 765 1324 769
rect 1328 765 1332 769
rect 1349 765 1353 769
rect 1357 765 1361 769
rect 1378 765 1382 769
rect 1812 765 1816 769
rect 1833 765 1837 769
rect 1841 765 1845 769
rect 1862 765 1866 769
rect 1870 765 1874 769
rect 1891 765 1895 769
rect 1899 765 1903 769
rect 1920 765 1924 769
rect 1928 765 1932 769
rect 1949 765 1953 769
rect 1957 765 1961 769
rect 1978 765 1982 769
rect 2415 768 2419 772
rect 2436 768 2440 772
rect 2444 768 2448 772
rect 2465 768 2469 772
rect 2473 768 2477 772
rect 2494 768 2498 772
rect 2502 768 2506 772
rect 2523 768 2527 772
rect 2531 768 2535 772
rect 2552 768 2556 772
rect 2560 768 2564 772
rect 2581 768 2585 772
rect -391 628 -386 633
rect -372 628 -367 633
rect -360 628 -355 633
rect -341 628 -336 633
rect -327 628 -322 633
rect -308 628 -303 633
rect -255 629 -250 634
rect -236 629 -231 634
rect -224 629 -219 634
rect -205 629 -200 634
rect -191 629 -186 634
rect -172 629 -167 634
rect -120 630 -115 635
rect -101 630 -96 635
rect -89 630 -84 635
rect -70 630 -65 635
rect -56 630 -51 635
rect -37 630 -32 635
rect 17 628 22 633
rect 36 628 41 633
rect 48 628 53 633
rect 67 628 72 633
rect 81 628 86 633
rect 100 628 105 633
rect -392 508 -387 513
rect -373 508 -368 513
rect -361 508 -356 513
rect -342 508 -337 513
rect -328 508 -323 513
rect -309 508 -304 513
rect -246 509 -241 514
rect -227 509 -222 514
rect -215 509 -210 514
rect -196 509 -191 514
rect -182 509 -177 514
rect -163 509 -158 514
rect -116 512 -111 517
rect -97 512 -92 517
rect -85 512 -80 517
rect -66 512 -61 517
rect -52 512 -47 517
rect -33 512 -28 517
rect 25 511 30 516
rect -1052 454 -1047 459
rect -1033 454 -1028 459
rect -1021 454 -1016 459
rect -1002 454 -997 459
rect -988 454 -983 459
rect -969 454 -964 459
rect 44 511 49 516
rect 56 511 61 516
rect 75 511 80 516
rect 89 511 94 516
rect 108 511 113 516
rect -1239 426 -1235 430
rect -1191 426 -1187 430
rect -1050 353 -1045 358
rect -1031 353 -1026 358
rect -1019 353 -1014 358
rect -1000 353 -995 358
rect -986 353 -981 358
rect -967 353 -962 358
rect -1047 254 -1042 259
rect -1028 254 -1023 259
rect -1016 254 -1011 259
rect -997 254 -992 259
rect -983 254 -978 259
rect -964 254 -959 259
rect -1241 207 -1237 211
rect -1193 207 -1189 211
rect -378 203 -373 208
rect -359 203 -354 208
rect -347 203 -342 208
rect -328 203 -323 208
rect -314 203 -309 208
rect -295 203 -290 208
rect -242 204 -237 209
rect -223 204 -218 209
rect -211 204 -206 209
rect -192 204 -187 209
rect -178 204 -173 209
rect -159 204 -154 209
rect -107 205 -102 210
rect -88 205 -83 210
rect -76 205 -71 210
rect -57 205 -52 210
rect -43 205 -38 210
rect -24 205 -19 210
rect 30 203 35 208
rect -1045 146 -1040 151
rect -1026 146 -1021 151
rect -1014 146 -1009 151
rect -995 146 -990 151
rect -981 146 -976 151
rect -962 146 -957 151
rect 49 203 54 208
rect 61 203 66 208
rect 80 203 85 208
rect 94 203 99 208
rect 113 203 118 208
rect -379 83 -374 88
rect -360 83 -355 88
rect -348 83 -343 88
rect -329 83 -324 88
rect -315 83 -310 88
rect -296 83 -291 88
rect -233 84 -228 89
rect -214 84 -209 89
rect -202 84 -197 89
rect -183 84 -178 89
rect -169 84 -164 89
rect -150 84 -145 89
rect -103 87 -98 92
rect -84 87 -79 92
rect -72 87 -67 92
rect -53 87 -48 92
rect -39 87 -34 92
rect -20 87 -15 92
rect 38 86 43 91
rect 57 86 62 91
rect 69 86 74 91
rect 88 86 93 91
rect 102 86 107 91
rect 121 86 126 91
rect 2077 10 2081 14
rect 2125 10 2129 14
rect 2602 11 2606 15
rect 2347 5 2351 9
rect 2395 5 2399 9
rect 2650 11 2654 15
rect 2870 11 2874 15
rect 2918 11 2922 15
rect 3426 -137 3430 -133
rect 3451 -137 3455 -133
rect 3460 -137 3464 -133
rect 3485 -137 3489 -133
rect 3493 -137 3497 -133
rect 3518 -137 3522 -133
rect 3526 -137 3530 -133
rect 3551 -137 3555 -133
rect 3559 -137 3563 -133
rect 3584 -137 3588 -133
rect 2219 -187 2223 -183
rect 2255 -187 2259 -183
rect 2263 -187 2267 -183
rect 2299 -187 2303 -183
rect 2307 -187 2311 -183
rect 2343 -187 2347 -183
rect 2351 -187 2355 -183
rect 2387 -187 2391 -183
rect 2395 -187 2399 -183
rect 2431 -187 2435 -183
rect 2439 -187 2443 -183
rect 2475 -187 2479 -183
rect 2601 -187 2605 -183
rect 2637 -187 2641 -183
rect 2645 -187 2649 -183
rect 2681 -187 2685 -183
rect 2689 -187 2693 -183
rect 2725 -187 2729 -183
rect 2733 -187 2737 -183
rect 2769 -187 2773 -183
rect 2777 -187 2781 -183
rect 2813 -187 2817 -183
rect 2821 -187 2825 -183
rect 2857 -187 2861 -183
rect 2983 -187 2987 -183
rect 3019 -187 3023 -183
rect 3027 -187 3031 -183
rect 3063 -187 3067 -183
rect 3071 -187 3075 -183
rect 3107 -187 3111 -183
rect 3115 -187 3119 -183
rect 3151 -187 3155 -183
rect 3159 -187 3163 -183
rect 3195 -187 3199 -183
rect 3203 -187 3207 -183
rect 3239 -187 3243 -183
rect -326 -247 -321 -242
rect -307 -247 -302 -242
rect -295 -247 -290 -242
rect -276 -247 -271 -242
rect -262 -247 -257 -242
rect -243 -247 -238 -242
rect -190 -246 -185 -241
rect -171 -246 -166 -241
rect -159 -246 -154 -241
rect -140 -246 -135 -241
rect -126 -246 -121 -241
rect -107 -246 -102 -241
rect -55 -245 -50 -240
rect -36 -245 -31 -240
rect -24 -245 -19 -240
rect -5 -245 0 -240
rect 9 -245 14 -240
rect 28 -245 33 -240
rect 82 -247 87 -242
rect 101 -247 106 -242
rect 113 -247 118 -242
rect 132 -247 137 -242
rect 146 -247 151 -242
rect 165 -247 170 -242
rect 2041 -259 2046 -254
rect 2060 -259 2065 -254
rect 2072 -259 2077 -254
rect 2091 -259 2096 -254
rect 2105 -259 2110 -254
rect 2124 -259 2129 -254
rect -327 -367 -322 -362
rect -308 -367 -303 -362
rect -296 -367 -291 -362
rect -277 -367 -272 -362
rect -263 -367 -258 -362
rect -244 -367 -239 -362
rect -181 -366 -176 -361
rect -162 -366 -157 -361
rect -150 -366 -145 -361
rect -131 -366 -126 -361
rect -117 -366 -112 -361
rect -98 -366 -93 -361
rect -51 -363 -46 -358
rect -32 -363 -27 -358
rect -20 -363 -15 -358
rect -1 -363 4 -358
rect 13 -363 18 -358
rect 32 -363 37 -358
rect 90 -364 95 -359
rect 109 -364 114 -359
rect 121 -364 126 -359
rect 140 -364 145 -359
rect 154 -364 159 -359
rect 173 -364 178 -359
rect 401 -427 406 -422
rect 420 -427 425 -422
rect 432 -427 437 -422
rect 451 -427 456 -422
rect 465 -427 470 -422
rect 484 -427 489 -422
rect 2057 -514 2061 -510
rect 2080 -514 2084 -510
rect 2091 -514 2095 -510
rect 2114 -514 2118 -510
rect 2124 -514 2128 -510
rect 2147 -514 2151 -510
rect 2156 -514 2160 -510
rect 2179 -514 2183 -510
rect 2188 -514 2192 -510
rect 2211 -514 2215 -510
rect 2220 -514 2224 -510
rect 2243 -514 2247 -510
rect -270 -533 -265 -528
rect -251 -533 -246 -528
rect -239 -533 -234 -528
rect -220 -533 -215 -528
rect -206 -533 -201 -528
rect -187 -533 -182 -528
rect -94 -589 -89 -584
rect -75 -589 -70 -584
rect -63 -589 -58 -584
rect -44 -589 -39 -584
rect -30 -589 -25 -584
rect -11 -589 -6 -584
rect 160 -599 165 -594
rect 179 -599 184 -594
rect 191 -599 196 -594
rect 210 -599 215 -594
rect 224 -599 229 -594
rect 243 -599 248 -594
rect 2056 -761 2060 -757
rect 2079 -761 2083 -757
rect 2090 -761 2094 -757
rect 2113 -761 2117 -757
rect 2123 -761 2127 -757
rect 2146 -761 2150 -757
rect 2155 -761 2159 -757
rect 2178 -761 2182 -757
rect 2187 -761 2191 -757
rect 2210 -761 2214 -757
rect 2219 -761 2223 -757
rect 2242 -761 2246 -757
rect 2410 -807 2414 -803
rect 2446 -807 2450 -803
rect 2454 -807 2458 -803
rect 2490 -807 2494 -803
rect 2498 -807 2502 -803
rect 2534 -807 2538 -803
rect 2542 -807 2546 -803
rect 2578 -807 2582 -803
rect 2586 -807 2590 -803
rect 2622 -807 2626 -803
rect 2630 -807 2634 -803
rect 2666 -807 2670 -803
rect 2060 -987 2064 -983
rect 2083 -987 2087 -983
rect 2094 -987 2098 -983
rect 2117 -987 2121 -983
rect 2127 -987 2131 -983
rect 2150 -987 2154 -983
rect 2159 -987 2163 -983
rect 2182 -987 2186 -983
rect 2191 -987 2195 -983
rect 2214 -987 2218 -983
rect 2223 -987 2227 -983
rect 2246 -987 2250 -983
rect 2057 -1194 2061 -1190
rect 2080 -1194 2084 -1190
rect 2091 -1194 2095 -1190
rect 2114 -1194 2118 -1190
rect 2124 -1194 2128 -1190
rect 2147 -1194 2151 -1190
rect 2156 -1194 2160 -1190
rect 2179 -1194 2183 -1190
rect 2188 -1194 2192 -1190
rect 2211 -1194 2215 -1190
rect 2220 -1194 2224 -1190
rect 2243 -1194 2247 -1190
rect 2084 -1404 2089 -1399
rect 2103 -1404 2108 -1399
rect 2115 -1404 2120 -1399
rect 2134 -1404 2139 -1399
rect 2148 -1404 2153 -1399
rect 2167 -1404 2172 -1399
rect 2270 -1413 2274 -1409
rect 2306 -1413 2310 -1409
rect 2314 -1413 2318 -1409
rect 2350 -1413 2354 -1409
rect 2358 -1413 2362 -1409
rect 2394 -1413 2398 -1409
rect 2402 -1413 2406 -1409
rect 2438 -1413 2442 -1409
rect 2446 -1413 2450 -1409
rect 2482 -1413 2486 -1409
rect 2490 -1413 2494 -1409
rect 2526 -1413 2530 -1409
rect 2642 -1412 2646 -1408
rect 2678 -1412 2682 -1408
rect 2686 -1412 2690 -1408
rect 2722 -1412 2726 -1408
rect 2730 -1412 2734 -1408
rect 2766 -1412 2770 -1408
rect 2774 -1412 2778 -1408
rect 2810 -1412 2814 -1408
rect 2818 -1412 2822 -1408
rect 2854 -1412 2858 -1408
rect 2862 -1412 2866 -1408
rect 2898 -1412 2902 -1408
rect 3016 -1412 3020 -1408
rect 3052 -1412 3056 -1408
rect 3060 -1412 3064 -1408
rect 3096 -1412 3100 -1408
rect 3104 -1412 3108 -1408
rect 3140 -1412 3144 -1408
rect 3148 -1412 3152 -1408
rect 3184 -1412 3188 -1408
rect 3192 -1412 3196 -1408
rect 3228 -1412 3232 -1408
rect 3236 -1412 3240 -1408
rect 3272 -1412 3276 -1408
rect 3476 -1464 3480 -1460
rect 3501 -1464 3505 -1460
rect 3510 -1464 3514 -1460
rect 3535 -1464 3539 -1460
rect 3543 -1464 3547 -1460
rect 3568 -1464 3572 -1460
rect 3576 -1464 3580 -1460
rect 3601 -1464 3605 -1460
rect 3609 -1464 3613 -1460
rect 3634 -1464 3638 -1460
rect 2104 -1529 2108 -1525
rect 2152 -1529 2156 -1525
rect 2301 -1575 2305 -1571
rect 2349 -1575 2353 -1571
rect 2709 -1599 2713 -1595
rect 2757 -1599 2761 -1595
rect 3136 -1598 3140 -1594
rect 3184 -1598 3188 -1594
<< polysilicon >>
rect 954 2049 1017 2051
rect 503 2047 566 2049
rect 503 2041 506 2047
rect 532 2041 534 2044
rect 563 2041 566 2047
rect 721 2047 784 2049
rect 592 2041 595 2045
rect 621 2041 624 2045
rect 651 2041 654 2045
rect 721 2041 724 2047
rect 750 2041 752 2044
rect 781 2041 784 2047
rect 810 2041 813 2045
rect 839 2041 842 2045
rect 869 2041 872 2045
rect 954 2043 957 2049
rect 983 2043 985 2046
rect 1014 2043 1017 2049
rect 1214 2050 1277 2052
rect 1043 2043 1046 2047
rect 1072 2043 1075 2047
rect 1102 2043 1105 2047
rect 1214 2044 1217 2050
rect 1243 2044 1245 2047
rect 1274 2044 1277 2050
rect 1303 2044 1306 2048
rect 1332 2044 1335 2048
rect 1362 2044 1365 2048
rect 503 1969 506 2034
rect 532 1969 534 2034
rect 563 1969 566 2034
rect 592 1969 595 2034
rect 614 2007 617 2012
rect 621 1969 624 2034
rect 651 1969 654 2034
rect 721 1969 724 2034
rect 750 1969 752 2034
rect 781 1969 784 2034
rect 810 1969 813 2034
rect 832 2007 835 2012
rect 839 1969 842 2034
rect 869 1969 872 2034
rect 954 1971 957 2036
rect 983 1971 985 2036
rect 1014 1971 1017 2036
rect 1043 1971 1046 2036
rect 1065 2009 1068 2014
rect 1072 1971 1075 2036
rect 1102 1971 1105 2036
rect 1214 1972 1217 2037
rect 1243 1972 1245 2037
rect 1274 1972 1277 2037
rect 1303 1972 1306 2037
rect 1325 2010 1328 2015
rect 1332 1972 1335 2037
rect 1362 1972 1365 2037
rect 503 1957 506 1962
rect 532 1950 534 1962
rect 563 1959 566 1962
rect 592 1950 595 1962
rect 621 1957 624 1962
rect 651 1957 654 1962
rect 721 1957 724 1962
rect 532 1948 595 1950
rect 750 1950 752 1962
rect 781 1959 784 1962
rect 810 1950 813 1962
rect 839 1957 842 1962
rect 869 1957 872 1962
rect 954 1959 957 1964
rect 750 1947 813 1950
rect 983 1952 985 1964
rect 1014 1961 1017 1964
rect 1043 1952 1046 1964
rect 1072 1959 1075 1964
rect 1102 1959 1105 1964
rect 1214 1960 1217 1965
rect 983 1949 1046 1952
rect 1243 1953 1245 1965
rect 1274 1962 1277 1965
rect 1303 1953 1306 1965
rect 1332 1960 1335 1965
rect 1362 1960 1365 1965
rect 1243 1950 1306 1953
rect 532 1849 595 1851
rect 2361 1849 2424 1851
rect 532 1843 535 1849
rect 561 1843 563 1846
rect 592 1843 595 1849
rect 621 1843 624 1847
rect 650 1843 653 1847
rect 680 1843 683 1847
rect 759 1843 763 1849
rect 791 1843 795 1847
rect 825 1843 829 1847
rect 1158 1846 1221 1848
rect 1758 1846 1821 1848
rect 532 1771 535 1836
rect 561 1771 563 1836
rect 592 1771 595 1836
rect 621 1771 624 1836
rect 643 1809 646 1814
rect 650 1771 653 1836
rect 680 1771 683 1836
rect 1158 1840 1161 1846
rect 1187 1840 1189 1843
rect 1218 1840 1221 1846
rect 1247 1840 1250 1844
rect 1276 1840 1279 1844
rect 1306 1840 1309 1844
rect 1385 1840 1389 1846
rect 1417 1840 1421 1844
rect 1451 1840 1455 1844
rect 1758 1840 1761 1846
rect 1787 1840 1789 1843
rect 1818 1840 1821 1846
rect 1847 1840 1850 1844
rect 1876 1840 1879 1844
rect 1906 1840 1909 1844
rect 1985 1840 1989 1846
rect 2017 1840 2021 1844
rect 2051 1840 2055 1844
rect 2361 1843 2364 1849
rect 2390 1843 2392 1846
rect 2421 1843 2424 1849
rect 2450 1843 2453 1847
rect 2479 1843 2482 1847
rect 2509 1843 2512 1847
rect 2588 1843 2592 1849
rect 2620 1843 2624 1847
rect 2654 1843 2658 1847
rect 759 1800 763 1834
rect 760 1795 763 1800
rect 759 1785 763 1795
rect 791 1785 795 1834
rect 825 1785 829 1834
rect 932 1818 934 1821
rect 950 1818 952 1821
rect 969 1818 971 1821
rect 932 1791 934 1814
rect 950 1793 952 1814
rect 969 1794 971 1814
rect 933 1787 934 1791
rect 951 1789 952 1793
rect 970 1790 971 1794
rect 932 1777 934 1787
rect 950 1777 952 1789
rect 969 1777 971 1790
rect 759 1773 763 1776
rect 791 1773 795 1776
rect 825 1773 829 1776
rect 932 1770 934 1773
rect 950 1770 952 1773
rect 969 1770 971 1773
rect 1158 1768 1161 1833
rect 1187 1768 1189 1833
rect 1218 1768 1221 1833
rect 1247 1768 1250 1833
rect 1269 1806 1272 1811
rect 1276 1768 1279 1833
rect 1306 1768 1309 1833
rect 1385 1797 1389 1831
rect 1386 1792 1389 1797
rect 1385 1782 1389 1792
rect 1417 1782 1421 1831
rect 1451 1782 1455 1831
rect 1558 1815 1560 1818
rect 1576 1815 1578 1818
rect 1595 1815 1597 1818
rect 1558 1788 1560 1811
rect 1576 1790 1578 1811
rect 1595 1791 1597 1811
rect 1559 1784 1560 1788
rect 1577 1786 1578 1790
rect 1596 1787 1597 1791
rect 1558 1774 1560 1784
rect 1576 1774 1578 1786
rect 1595 1774 1597 1787
rect 1385 1770 1389 1773
rect 1417 1770 1421 1773
rect 1451 1770 1455 1773
rect 532 1759 535 1764
rect 561 1752 563 1764
rect 592 1761 595 1764
rect 621 1752 624 1764
rect 650 1759 653 1764
rect 680 1759 683 1764
rect 1558 1767 1560 1770
rect 1576 1767 1578 1770
rect 1595 1767 1597 1770
rect 1758 1768 1761 1833
rect 1787 1768 1789 1833
rect 1818 1768 1821 1833
rect 1847 1768 1850 1833
rect 1869 1806 1872 1811
rect 1876 1768 1879 1833
rect 1906 1768 1909 1833
rect 1985 1797 1989 1831
rect 1986 1792 1989 1797
rect 1985 1782 1989 1792
rect 2017 1782 2021 1831
rect 2051 1782 2055 1831
rect 2158 1815 2160 1818
rect 2176 1815 2178 1818
rect 2195 1815 2197 1818
rect 2158 1788 2160 1811
rect 2176 1790 2178 1811
rect 2195 1791 2197 1811
rect 2159 1784 2160 1788
rect 2177 1786 2178 1790
rect 2196 1787 2197 1791
rect 2158 1774 2160 1784
rect 2176 1774 2178 1786
rect 2195 1774 2197 1787
rect 1985 1770 1989 1773
rect 2017 1770 2021 1773
rect 2051 1770 2055 1773
rect 2361 1771 2364 1836
rect 2390 1771 2392 1836
rect 2421 1771 2424 1836
rect 2450 1771 2453 1836
rect 2472 1809 2475 1814
rect 2479 1771 2482 1836
rect 2509 1771 2512 1836
rect 2588 1800 2592 1834
rect 2589 1795 2592 1800
rect 2588 1785 2592 1795
rect 2620 1785 2624 1834
rect 2654 1785 2658 1834
rect 2761 1818 2763 1821
rect 2779 1818 2781 1821
rect 2798 1818 2800 1821
rect 2761 1791 2763 1814
rect 2779 1793 2781 1814
rect 2798 1794 2800 1814
rect 2762 1787 2763 1791
rect 2780 1789 2781 1793
rect 2799 1790 2800 1794
rect 2761 1777 2763 1787
rect 2779 1777 2781 1789
rect 2798 1777 2800 1790
rect 2588 1773 2592 1776
rect 2620 1773 2624 1776
rect 2654 1773 2658 1776
rect 2158 1767 2160 1770
rect 2176 1767 2178 1770
rect 2195 1767 2197 1770
rect 2761 1770 2763 1773
rect 2779 1770 2781 1773
rect 2798 1770 2800 1773
rect 1158 1756 1161 1761
rect 561 1749 624 1752
rect 1187 1749 1189 1761
rect 1218 1758 1221 1761
rect 1247 1749 1250 1761
rect 1276 1756 1279 1761
rect 1306 1756 1309 1761
rect 1758 1756 1761 1761
rect 1187 1746 1250 1749
rect 1787 1749 1789 1761
rect 1818 1758 1821 1761
rect 1847 1749 1850 1761
rect 1876 1756 1879 1761
rect 1906 1756 1909 1761
rect 2361 1759 2364 1764
rect 2390 1752 2392 1764
rect 2421 1761 2424 1764
rect 2450 1752 2453 1764
rect 2479 1759 2482 1764
rect 2509 1759 2512 1764
rect 2390 1749 2453 1752
rect 1787 1746 1850 1749
rect 775 1704 779 1710
rect 807 1704 811 1708
rect 841 1704 845 1708
rect 1401 1701 1405 1707
rect 1433 1701 1437 1705
rect 1467 1701 1471 1705
rect 2001 1701 2005 1707
rect 2033 1701 2037 1705
rect 2067 1701 2071 1705
rect 2604 1704 2608 1710
rect 2636 1704 2640 1708
rect 2670 1704 2674 1708
rect 775 1661 779 1695
rect 776 1656 779 1661
rect 775 1646 779 1656
rect 807 1646 811 1695
rect 841 1646 845 1695
rect 1401 1658 1405 1692
rect 1402 1653 1405 1658
rect 1401 1643 1405 1653
rect 1433 1643 1437 1692
rect 1467 1643 1471 1692
rect 2001 1658 2005 1692
rect 2002 1653 2005 1658
rect 2001 1643 2005 1653
rect 2033 1643 2037 1692
rect 2067 1643 2071 1692
rect 2604 1661 2608 1695
rect 2605 1656 2608 1661
rect 2604 1646 2608 1656
rect 2636 1646 2640 1695
rect 2670 1646 2674 1695
rect 775 1634 779 1637
rect 807 1634 811 1637
rect 841 1634 845 1637
rect 2604 1634 2608 1637
rect 2636 1634 2640 1637
rect 2670 1634 2674 1637
rect 1401 1631 1405 1634
rect 1433 1631 1437 1634
rect 1467 1631 1471 1634
rect 2001 1631 2005 1634
rect 2033 1631 2037 1634
rect 2067 1631 2071 1634
rect 542 1593 605 1595
rect 542 1587 545 1593
rect 571 1587 573 1590
rect 602 1587 605 1593
rect 2371 1593 2434 1595
rect 631 1587 634 1591
rect 660 1587 663 1591
rect 690 1587 693 1591
rect 1168 1590 1231 1592
rect 1168 1584 1171 1590
rect 1197 1584 1199 1587
rect 1228 1584 1231 1590
rect 1768 1590 1831 1592
rect 1257 1584 1260 1588
rect 1286 1584 1289 1588
rect 1316 1584 1319 1588
rect 1768 1584 1771 1590
rect 1797 1584 1799 1587
rect 1828 1584 1831 1590
rect 1857 1584 1860 1588
rect 1886 1584 1889 1588
rect 1916 1584 1919 1588
rect 2371 1587 2374 1593
rect 2400 1587 2402 1590
rect 2431 1587 2434 1593
rect 2460 1587 2463 1591
rect 2489 1587 2492 1591
rect 2519 1587 2522 1591
rect 542 1515 545 1580
rect 571 1515 573 1580
rect 602 1515 605 1580
rect 631 1515 634 1580
rect 653 1553 656 1558
rect 660 1515 663 1580
rect 690 1515 693 1580
rect 1168 1512 1171 1577
rect 1197 1512 1199 1577
rect 1228 1512 1231 1577
rect 1257 1512 1260 1577
rect 1279 1550 1282 1555
rect 1286 1512 1289 1577
rect 1316 1512 1319 1577
rect 1768 1512 1771 1577
rect 1797 1512 1799 1577
rect 1828 1512 1831 1577
rect 1857 1512 1860 1577
rect 1879 1550 1882 1555
rect 1886 1512 1889 1577
rect 1916 1512 1919 1577
rect 2371 1515 2374 1580
rect 2400 1515 2402 1580
rect 2431 1515 2434 1580
rect 2460 1515 2463 1580
rect 2482 1553 2485 1558
rect 2489 1515 2492 1580
rect 2519 1515 2522 1580
rect 542 1503 545 1508
rect 571 1496 573 1508
rect 602 1505 605 1508
rect 631 1496 634 1508
rect 660 1503 663 1508
rect 690 1503 693 1508
rect 1168 1500 1171 1505
rect 571 1493 634 1496
rect 1197 1493 1199 1505
rect 1228 1502 1231 1505
rect 1257 1493 1260 1505
rect 1286 1500 1289 1505
rect 1316 1500 1319 1505
rect 1768 1500 1771 1505
rect 1197 1490 1260 1493
rect 1797 1493 1799 1505
rect 1828 1502 1831 1505
rect 1857 1493 1860 1505
rect 1886 1500 1889 1505
rect 1916 1500 1919 1505
rect 2371 1503 2374 1508
rect 2400 1496 2402 1508
rect 2431 1505 2434 1508
rect 2460 1496 2463 1508
rect 2489 1503 2492 1508
rect 2519 1503 2522 1508
rect 2400 1493 2463 1496
rect 1797 1490 1860 1493
rect 1007 1234 1070 1236
rect 556 1232 619 1234
rect 556 1226 559 1232
rect 585 1226 587 1229
rect 616 1226 619 1232
rect 774 1232 837 1234
rect 645 1226 648 1230
rect 674 1226 677 1230
rect 704 1226 707 1230
rect 774 1226 777 1232
rect 803 1226 805 1229
rect 834 1226 837 1232
rect 863 1226 866 1230
rect 892 1226 895 1230
rect 922 1226 925 1230
rect 1007 1228 1010 1234
rect 1036 1228 1038 1231
rect 1067 1228 1070 1234
rect 1267 1235 1330 1237
rect 1096 1228 1099 1232
rect 1125 1228 1128 1232
rect 1155 1228 1158 1232
rect 1267 1229 1270 1235
rect 1296 1229 1298 1232
rect 1327 1229 1330 1235
rect 1356 1229 1359 1233
rect 1385 1229 1388 1233
rect 1415 1229 1418 1233
rect 556 1154 559 1219
rect 585 1154 587 1219
rect 616 1154 619 1219
rect 645 1154 648 1219
rect 667 1192 670 1197
rect 674 1154 677 1219
rect 704 1154 707 1219
rect 774 1154 777 1219
rect 803 1154 805 1219
rect 834 1154 837 1219
rect 863 1154 866 1219
rect 885 1192 888 1197
rect 892 1154 895 1219
rect 922 1154 925 1219
rect 1007 1156 1010 1221
rect 1036 1156 1038 1221
rect 1067 1156 1070 1221
rect 1096 1156 1099 1221
rect 1118 1194 1121 1199
rect 1125 1156 1128 1221
rect 1155 1156 1158 1221
rect 1267 1157 1270 1222
rect 1296 1157 1298 1222
rect 1327 1157 1330 1222
rect 1356 1157 1359 1222
rect 1378 1195 1381 1200
rect 1385 1157 1388 1222
rect 1415 1157 1418 1222
rect 556 1142 559 1147
rect 585 1135 587 1147
rect 616 1144 619 1147
rect 645 1135 648 1147
rect 674 1142 677 1147
rect 704 1142 707 1147
rect 774 1142 777 1147
rect 585 1133 648 1135
rect 803 1135 805 1147
rect 834 1144 837 1147
rect 863 1135 866 1147
rect 892 1142 895 1147
rect 922 1142 925 1147
rect 1007 1144 1010 1149
rect 803 1132 866 1135
rect 1036 1137 1038 1149
rect 1067 1146 1070 1149
rect 1096 1137 1099 1149
rect 1125 1144 1128 1149
rect 1155 1144 1158 1149
rect 1267 1145 1270 1150
rect 1036 1134 1099 1137
rect 1296 1138 1298 1150
rect 1327 1147 1330 1150
rect 1356 1138 1359 1150
rect 1385 1145 1388 1150
rect 1415 1145 1418 1150
rect 1296 1135 1359 1138
rect -401 1076 -397 1082
rect -369 1076 -365 1080
rect -335 1076 -331 1080
rect -265 1077 -261 1083
rect -233 1077 -229 1081
rect -199 1077 -195 1081
rect -130 1078 -126 1084
rect -98 1078 -94 1082
rect -64 1078 -60 1082
rect 7 1076 11 1082
rect 39 1076 43 1080
rect 73 1076 77 1080
rect -401 1033 -397 1067
rect -400 1028 -397 1033
rect -401 1018 -397 1028
rect -369 1018 -365 1067
rect -335 1018 -331 1067
rect -265 1034 -261 1068
rect -264 1029 -261 1034
rect -265 1019 -261 1029
rect -233 1019 -229 1068
rect -199 1019 -195 1068
rect -130 1035 -126 1069
rect -129 1030 -126 1035
rect -130 1020 -126 1030
rect -98 1020 -94 1069
rect -64 1020 -60 1069
rect 7 1033 11 1067
rect 8 1028 11 1033
rect 7 1018 11 1028
rect 39 1018 43 1067
rect 73 1018 77 1067
rect 585 1034 648 1036
rect 2414 1034 2477 1036
rect 585 1028 588 1034
rect 614 1028 616 1031
rect 645 1028 648 1034
rect 674 1028 677 1032
rect 703 1028 706 1032
rect 733 1028 736 1032
rect 812 1028 816 1034
rect 844 1028 848 1032
rect 878 1028 882 1032
rect 1211 1031 1274 1033
rect 1811 1031 1874 1033
rect -401 1006 -397 1009
rect -369 1006 -365 1009
rect -335 1006 -331 1009
rect -265 1007 -261 1010
rect -233 1007 -229 1010
rect -199 1007 -195 1010
rect -130 1008 -126 1011
rect -98 1008 -94 1011
rect -64 1008 -60 1011
rect 7 1006 11 1009
rect 39 1006 43 1009
rect 73 1006 77 1009
rect -402 956 -398 962
rect -370 956 -366 960
rect -336 956 -332 960
rect -256 957 -252 963
rect -224 957 -220 961
rect -190 957 -186 961
rect -126 960 -122 966
rect -94 960 -90 964
rect -60 960 -56 964
rect 15 959 19 965
rect 47 959 51 963
rect 81 959 85 963
rect -402 913 -398 947
rect -401 908 -398 913
rect -402 898 -398 908
rect -370 898 -366 947
rect -336 898 -332 947
rect -256 914 -252 948
rect -255 909 -252 914
rect -256 899 -252 909
rect -224 899 -220 948
rect -190 899 -186 948
rect -126 917 -122 951
rect -125 912 -122 917
rect -126 902 -122 912
rect -94 902 -90 951
rect -60 902 -56 951
rect 585 956 588 1021
rect 614 956 616 1021
rect 645 956 648 1021
rect 674 956 677 1021
rect 696 994 699 999
rect 703 956 706 1021
rect 733 956 736 1021
rect 1211 1025 1214 1031
rect 1240 1025 1242 1028
rect 1271 1025 1274 1031
rect 1300 1025 1303 1029
rect 1329 1025 1332 1029
rect 1359 1025 1362 1029
rect 1438 1025 1442 1031
rect 1470 1025 1474 1029
rect 1504 1025 1508 1029
rect 1811 1025 1814 1031
rect 1840 1025 1842 1028
rect 1871 1025 1874 1031
rect 1900 1025 1903 1029
rect 1929 1025 1932 1029
rect 1959 1025 1962 1029
rect 2038 1025 2042 1031
rect 2070 1025 2074 1029
rect 2104 1025 2108 1029
rect 2414 1028 2417 1034
rect 2443 1028 2445 1031
rect 2474 1028 2477 1034
rect 2503 1028 2506 1032
rect 2532 1028 2535 1032
rect 2562 1028 2565 1032
rect 2641 1028 2645 1034
rect 2673 1028 2677 1032
rect 2707 1028 2711 1032
rect 812 985 816 1019
rect 813 980 816 985
rect 812 970 816 980
rect 844 970 848 1019
rect 878 970 882 1019
rect 985 1003 987 1006
rect 1003 1003 1005 1006
rect 1022 1003 1024 1006
rect 985 976 987 999
rect 1003 978 1005 999
rect 1022 979 1024 999
rect 986 972 987 976
rect 1004 974 1005 978
rect 1023 975 1024 979
rect 985 962 987 972
rect 1003 962 1005 974
rect 1022 962 1024 975
rect 812 958 816 961
rect 844 958 848 961
rect 878 958 882 961
rect 15 916 19 950
rect 16 911 19 916
rect 15 901 19 911
rect 47 901 51 950
rect 81 901 85 950
rect 985 955 987 958
rect 1003 955 1005 958
rect 1022 955 1024 958
rect 1211 953 1214 1018
rect 1240 953 1242 1018
rect 1271 953 1274 1018
rect 1300 953 1303 1018
rect 1322 991 1325 996
rect 1329 953 1332 1018
rect 1359 953 1362 1018
rect 1438 982 1442 1016
rect 1439 977 1442 982
rect 1438 967 1442 977
rect 1470 967 1474 1016
rect 1504 967 1508 1016
rect 1611 1000 1613 1003
rect 1629 1000 1631 1003
rect 1648 1000 1650 1003
rect 1611 973 1613 996
rect 1629 975 1631 996
rect 1648 976 1650 996
rect 1612 969 1613 973
rect 1630 971 1631 975
rect 1649 972 1650 976
rect 1611 959 1613 969
rect 1629 959 1631 971
rect 1648 959 1650 972
rect 1438 955 1442 958
rect 1470 955 1474 958
rect 1504 955 1508 958
rect 585 944 588 949
rect 614 937 616 949
rect 645 946 648 949
rect 674 937 677 949
rect 703 944 706 949
rect 733 944 736 949
rect 1611 952 1613 955
rect 1629 952 1631 955
rect 1648 952 1650 955
rect 1811 953 1814 1018
rect 1840 953 1842 1018
rect 1871 953 1874 1018
rect 1900 953 1903 1018
rect 1922 991 1925 996
rect 1929 953 1932 1018
rect 1959 953 1962 1018
rect 2038 982 2042 1016
rect 2039 977 2042 982
rect 2038 967 2042 977
rect 2070 967 2074 1016
rect 2104 967 2108 1016
rect 2211 1000 2213 1003
rect 2229 1000 2231 1003
rect 2248 1000 2250 1003
rect 2211 973 2213 996
rect 2229 975 2231 996
rect 2248 976 2250 996
rect 2212 969 2213 973
rect 2230 971 2231 975
rect 2249 972 2250 976
rect 2211 959 2213 969
rect 2229 959 2231 971
rect 2248 959 2250 972
rect 2038 955 2042 958
rect 2070 955 2074 958
rect 2104 955 2108 958
rect 2414 956 2417 1021
rect 2443 956 2445 1021
rect 2474 956 2477 1021
rect 2503 956 2506 1021
rect 2525 994 2528 999
rect 2532 956 2535 1021
rect 2562 956 2565 1021
rect 2641 985 2645 1019
rect 2642 980 2645 985
rect 2641 970 2645 980
rect 2673 970 2677 1019
rect 2707 970 2711 1019
rect 2814 1003 2816 1006
rect 2832 1003 2834 1006
rect 2851 1003 2853 1006
rect 2814 976 2816 999
rect 2832 978 2834 999
rect 2851 979 2853 999
rect 2815 972 2816 976
rect 2833 974 2834 978
rect 2852 975 2853 979
rect 2814 962 2816 972
rect 2832 962 2834 974
rect 2851 962 2853 975
rect 2641 958 2645 961
rect 2673 958 2677 961
rect 2707 958 2711 961
rect 2211 952 2213 955
rect 2229 952 2231 955
rect 2248 952 2250 955
rect 2814 955 2816 958
rect 2832 955 2834 958
rect 2851 955 2853 958
rect 1211 941 1214 946
rect 614 934 677 937
rect 1240 934 1242 946
rect 1271 943 1274 946
rect 1300 934 1303 946
rect 1329 941 1332 946
rect 1359 941 1362 946
rect 1811 941 1814 946
rect 1240 931 1303 934
rect 1840 934 1842 946
rect 1871 943 1874 946
rect 1900 934 1903 946
rect 1929 941 1932 946
rect 1959 941 1962 946
rect 2414 944 2417 949
rect 2443 937 2445 949
rect 2474 946 2477 949
rect 2503 937 2506 949
rect 2532 944 2535 949
rect 2562 944 2565 949
rect 2443 934 2506 937
rect 1840 931 1903 934
rect -126 890 -122 893
rect -94 890 -90 893
rect -60 890 -56 893
rect -402 886 -398 889
rect -370 886 -366 889
rect -336 886 -332 889
rect -256 887 -252 890
rect -224 887 -220 890
rect -190 887 -186 890
rect 15 889 19 892
rect 47 889 51 892
rect 81 889 85 892
rect 828 889 832 895
rect 860 889 864 893
rect 894 889 898 893
rect 1454 886 1458 892
rect 1486 886 1490 890
rect 1520 886 1524 890
rect 2054 886 2058 892
rect 2086 886 2090 890
rect 2120 886 2124 890
rect 2657 889 2661 895
rect 2689 889 2693 893
rect 2723 889 2727 893
rect 828 846 832 880
rect 829 841 832 846
rect 828 831 832 841
rect 860 831 864 880
rect 894 831 898 880
rect 1454 843 1458 877
rect 1455 838 1458 843
rect 1454 828 1458 838
rect 1486 828 1490 877
rect 1520 828 1524 877
rect 2054 843 2058 877
rect 2055 838 2058 843
rect 2054 828 2058 838
rect 2086 828 2090 877
rect 2120 828 2124 877
rect 2657 846 2661 880
rect 2658 841 2661 846
rect 2657 831 2661 841
rect 2689 831 2693 880
rect 2723 831 2727 880
rect 828 819 832 822
rect 860 819 864 822
rect 894 819 898 822
rect 2657 819 2661 822
rect 2689 819 2693 822
rect 2723 819 2727 822
rect 1454 816 1458 819
rect 1486 816 1490 819
rect 1520 816 1524 819
rect 2054 816 2058 819
rect 2086 816 2090 819
rect 2120 816 2124 819
rect 595 778 658 780
rect 595 772 598 778
rect 624 772 626 775
rect 655 772 658 778
rect 2424 778 2487 780
rect 684 772 687 776
rect 713 772 716 776
rect 743 772 746 776
rect 1221 775 1284 777
rect 1221 769 1224 775
rect 1250 769 1252 772
rect 1281 769 1284 775
rect 1821 775 1884 777
rect 1310 769 1313 773
rect 1339 769 1342 773
rect 1369 769 1372 773
rect 1821 769 1824 775
rect 1850 769 1852 772
rect 1881 769 1884 775
rect 1910 769 1913 773
rect 1939 769 1942 773
rect 1969 769 1972 773
rect 2424 772 2427 778
rect 2453 772 2455 775
rect 2484 772 2487 778
rect 2513 772 2516 776
rect 2542 772 2545 776
rect 2572 772 2575 776
rect 595 700 598 765
rect 624 700 626 765
rect 655 700 658 765
rect 684 700 687 765
rect 706 738 709 743
rect 713 700 716 765
rect 743 700 746 765
rect 1221 697 1224 762
rect 1250 697 1252 762
rect 1281 697 1284 762
rect 1310 697 1313 762
rect 1332 735 1335 740
rect 1339 697 1342 762
rect 1369 697 1372 762
rect 1821 697 1824 762
rect 1850 697 1852 762
rect 1881 697 1884 762
rect 1910 697 1913 762
rect 1932 735 1935 740
rect 1939 697 1942 762
rect 1969 697 1972 762
rect 2424 700 2427 765
rect 2453 700 2455 765
rect 2484 700 2487 765
rect 2513 700 2516 765
rect 2535 738 2538 743
rect 2542 700 2545 765
rect 2572 700 2575 765
rect 595 688 598 693
rect 624 681 626 693
rect 655 690 658 693
rect 684 681 687 693
rect 713 688 716 693
rect 743 688 746 693
rect 1221 685 1224 690
rect 624 678 687 681
rect 1250 678 1252 690
rect 1281 687 1284 690
rect 1310 678 1313 690
rect 1339 685 1342 690
rect 1369 685 1372 690
rect 1821 685 1824 690
rect 1250 675 1313 678
rect 1850 678 1852 690
rect 1881 687 1884 690
rect 1910 678 1913 690
rect 1939 685 1942 690
rect 1969 685 1972 690
rect 2424 688 2427 693
rect 2453 681 2455 693
rect 2484 690 2487 693
rect 2513 681 2516 693
rect 2542 688 2545 693
rect 2572 688 2575 693
rect 2453 678 2516 681
rect 1850 675 1913 678
rect -382 633 -378 639
rect -350 633 -346 637
rect -316 633 -312 637
rect -246 634 -242 640
rect -214 634 -210 638
rect -180 634 -176 638
rect -111 635 -107 641
rect -79 635 -75 639
rect -45 635 -41 639
rect 26 633 30 639
rect 58 633 62 637
rect 92 633 96 637
rect -382 590 -378 624
rect -381 585 -378 590
rect -382 575 -378 585
rect -350 575 -346 624
rect -316 575 -312 624
rect -246 591 -242 625
rect -245 586 -242 591
rect -246 576 -242 586
rect -214 576 -210 625
rect -180 576 -176 625
rect -111 592 -107 626
rect -110 587 -107 592
rect -111 577 -107 587
rect -79 577 -75 626
rect -45 577 -41 626
rect 26 590 30 624
rect 27 585 30 590
rect 26 575 30 585
rect 58 575 62 624
rect 92 575 96 624
rect -382 563 -378 566
rect -350 563 -346 566
rect -316 563 -312 566
rect -246 564 -242 567
rect -214 564 -210 567
rect -180 564 -176 567
rect -111 565 -107 568
rect -79 565 -75 568
rect -45 565 -41 568
rect 26 563 30 566
rect 58 563 62 566
rect 92 563 96 566
rect -383 513 -379 519
rect -351 513 -347 517
rect -317 513 -313 517
rect -237 514 -233 520
rect -205 514 -201 518
rect -171 514 -167 518
rect -107 517 -103 523
rect -75 517 -71 521
rect -41 517 -37 521
rect 34 516 38 522
rect 66 516 70 520
rect 100 516 104 520
rect -383 470 -379 504
rect -382 465 -379 470
rect -1043 459 -1039 465
rect -1011 459 -1007 463
rect -977 459 -973 463
rect -383 455 -379 465
rect -351 455 -347 504
rect -317 455 -313 504
rect -237 471 -233 505
rect -236 466 -233 471
rect -237 456 -233 466
rect -205 456 -201 505
rect -171 456 -167 505
rect -107 474 -103 508
rect -106 469 -103 474
rect -107 459 -103 469
rect -75 459 -71 508
rect -41 459 -37 508
rect 34 473 38 507
rect 35 468 38 473
rect -1215 430 -1211 442
rect -1215 392 -1211 420
rect -1043 416 -1039 450
rect -1042 411 -1039 416
rect -1043 401 -1039 411
rect -1011 401 -1007 450
rect -977 401 -973 450
rect 34 458 38 468
rect 66 458 70 507
rect 100 458 104 507
rect -107 447 -103 450
rect -75 447 -71 450
rect -41 447 -37 450
rect -383 443 -379 446
rect -351 443 -347 446
rect -317 443 -313 446
rect -237 444 -233 447
rect -205 444 -201 447
rect -171 444 -167 447
rect 34 446 38 449
rect 66 446 70 449
rect 100 446 104 449
rect -1043 389 -1039 392
rect -1011 389 -1007 392
rect -977 389 -973 392
rect -1215 363 -1211 378
rect -1041 358 -1037 364
rect -1009 358 -1005 362
rect -975 358 -971 362
rect -1041 315 -1037 349
rect -1040 310 -1037 315
rect -1041 300 -1037 310
rect -1009 300 -1005 349
rect -975 300 -971 349
rect -1041 288 -1037 291
rect -1009 288 -1005 291
rect -975 288 -971 291
rect -1038 259 -1034 265
rect -1006 259 -1002 263
rect -972 259 -968 263
rect -1217 211 -1213 223
rect -1038 216 -1034 250
rect -1037 211 -1034 216
rect -1038 201 -1034 211
rect -1006 201 -1002 250
rect -972 201 -968 250
rect -369 208 -365 214
rect -337 208 -333 212
rect -303 208 -299 212
rect -233 209 -229 215
rect -201 209 -197 213
rect -167 209 -163 213
rect -98 210 -94 216
rect -66 210 -62 214
rect -32 210 -28 214
rect -1217 173 -1213 201
rect 39 208 43 214
rect 71 208 75 212
rect 105 208 109 212
rect -1038 189 -1034 192
rect -1006 189 -1002 192
rect -972 189 -968 192
rect -369 165 -365 199
rect -368 160 -365 165
rect -1217 144 -1213 159
rect -1036 151 -1032 157
rect -1004 151 -1000 155
rect -970 151 -966 155
rect -369 150 -365 160
rect -337 150 -333 199
rect -303 150 -299 199
rect -233 166 -229 200
rect -232 161 -229 166
rect -233 151 -229 161
rect -201 151 -197 200
rect -167 151 -163 200
rect -98 167 -94 201
rect -97 162 -94 167
rect -98 152 -94 162
rect -66 152 -62 201
rect -32 152 -28 201
rect 39 165 43 199
rect 40 160 43 165
rect -1036 108 -1032 142
rect -1035 103 -1032 108
rect -1036 93 -1032 103
rect -1004 93 -1000 142
rect -970 93 -966 142
rect 39 150 43 160
rect 71 150 75 199
rect 105 150 109 199
rect -369 138 -365 141
rect -337 138 -333 141
rect -303 138 -299 141
rect -233 139 -229 142
rect -201 139 -197 142
rect -167 139 -163 142
rect -98 140 -94 143
rect -66 140 -62 143
rect -32 140 -28 143
rect 39 138 43 141
rect 71 138 75 141
rect 105 138 109 141
rect -370 88 -366 94
rect -338 88 -334 92
rect -304 88 -300 92
rect -224 89 -220 95
rect -192 89 -188 93
rect -158 89 -154 93
rect -94 92 -90 98
rect -62 92 -58 96
rect -28 92 -24 96
rect -1036 81 -1032 84
rect -1004 81 -1000 84
rect -970 81 -966 84
rect 47 91 51 97
rect 79 91 83 95
rect 113 91 117 95
rect -370 45 -366 79
rect -369 40 -366 45
rect -370 30 -366 40
rect -338 30 -334 79
rect -304 30 -300 79
rect -224 46 -220 80
rect -223 41 -220 46
rect -224 31 -220 41
rect -192 31 -188 80
rect -158 31 -154 80
rect -94 49 -90 83
rect -93 44 -90 49
rect -94 34 -90 44
rect -62 34 -58 83
rect -28 34 -24 83
rect 47 48 51 82
rect 48 43 51 48
rect 47 33 51 43
rect 79 33 83 82
rect 113 33 117 82
rect -94 22 -90 25
rect -62 22 -58 25
rect -28 22 -24 25
rect -370 18 -366 21
rect -338 18 -334 21
rect -304 18 -300 21
rect -224 19 -220 22
rect -192 19 -188 22
rect -158 19 -154 22
rect 47 21 51 24
rect 79 21 83 24
rect 113 21 117 24
rect 2101 14 2105 26
rect 2371 9 2375 21
rect 2626 15 2630 27
rect 2894 15 2898 27
rect 2101 -24 2105 4
rect 2371 -29 2375 -1
rect 2626 -23 2630 5
rect 2894 -23 2898 5
rect 2101 -53 2105 -38
rect 2371 -58 2375 -43
rect 2626 -52 2630 -37
rect 2894 -52 2898 -37
rect 3438 -133 3442 -123
rect 3473 -133 3477 -123
rect 3506 -133 3510 -123
rect 3539 -133 3543 -123
rect 3572 -133 3576 -123
rect 2235 -183 2239 -178
rect 2281 -183 2285 -178
rect 2326 -183 2330 -178
rect 2369 -183 2373 -178
rect 2414 -183 2418 -178
rect 2457 -183 2461 -178
rect 2617 -183 2621 -178
rect 2663 -183 2667 -178
rect 2708 -183 2712 -178
rect 2751 -183 2755 -178
rect 2796 -183 2800 -178
rect 2839 -183 2843 -178
rect 2999 -183 3003 -178
rect 3045 -183 3049 -178
rect 3090 -183 3094 -178
rect 3133 -183 3137 -178
rect 3178 -183 3182 -178
rect 3221 -183 3225 -178
rect -317 -242 -313 -236
rect -285 -242 -281 -238
rect -251 -242 -247 -238
rect -181 -241 -177 -235
rect -149 -241 -145 -237
rect -115 -241 -111 -237
rect -46 -240 -42 -234
rect -14 -240 -10 -236
rect 20 -240 24 -236
rect 91 -242 95 -236
rect 123 -242 127 -238
rect 157 -242 161 -238
rect -317 -285 -313 -251
rect -316 -290 -313 -285
rect -317 -300 -313 -290
rect -285 -300 -281 -251
rect -251 -300 -247 -251
rect -181 -284 -177 -250
rect -180 -289 -177 -284
rect -181 -299 -177 -289
rect -149 -299 -145 -250
rect -115 -299 -111 -250
rect -46 -283 -42 -249
rect -45 -288 -42 -283
rect -46 -298 -42 -288
rect -14 -298 -10 -249
rect 20 -298 24 -249
rect 91 -285 95 -251
rect 92 -290 95 -285
rect 91 -300 95 -290
rect 123 -300 127 -251
rect 157 -300 161 -251
rect 2050 -254 2054 -248
rect 2082 -254 2086 -250
rect 2116 -254 2120 -250
rect 2050 -297 2054 -263
rect -317 -312 -313 -309
rect -285 -312 -281 -309
rect -251 -312 -247 -309
rect -181 -311 -177 -308
rect -149 -311 -145 -308
rect -115 -311 -111 -308
rect -46 -310 -42 -307
rect -14 -310 -10 -307
rect 20 -310 24 -307
rect 2051 -302 2054 -297
rect 91 -312 95 -309
rect 123 -312 127 -309
rect 157 -312 161 -309
rect 2050 -312 2054 -302
rect 2082 -312 2086 -263
rect 2116 -312 2120 -263
rect 2235 -286 2239 -194
rect 2281 -241 2285 -194
rect 2280 -250 2285 -241
rect 2326 -242 2330 -194
rect 2369 -242 2373 -194
rect 2281 -286 2285 -250
rect 2328 -251 2330 -242
rect 2371 -251 2373 -242
rect 2414 -244 2418 -194
rect 2326 -286 2330 -251
rect 2369 -286 2373 -251
rect 2415 -253 2418 -244
rect 2414 -286 2418 -253
rect 2457 -286 2461 -194
rect 2617 -286 2621 -194
rect 2663 -241 2667 -194
rect 2662 -250 2667 -241
rect 2708 -242 2712 -194
rect 2751 -242 2755 -194
rect 2663 -286 2667 -250
rect 2710 -251 2712 -242
rect 2753 -251 2755 -242
rect 2796 -244 2800 -194
rect 2708 -286 2712 -251
rect 2751 -286 2755 -251
rect 2797 -253 2800 -244
rect 2796 -286 2800 -253
rect 2839 -286 2843 -194
rect 2999 -286 3003 -194
rect 3045 -241 3049 -194
rect 3044 -250 3049 -241
rect 3090 -242 3094 -194
rect 3133 -242 3137 -194
rect 3045 -286 3049 -250
rect 3092 -251 3094 -242
rect 3135 -251 3137 -242
rect 3178 -244 3182 -194
rect 3090 -286 3094 -251
rect 3133 -286 3137 -251
rect 3179 -253 3182 -244
rect 3178 -286 3182 -253
rect 3221 -286 3225 -194
rect 3438 -215 3442 -142
rect 3473 -215 3477 -142
rect 3506 -215 3510 -142
rect 3539 -215 3543 -142
rect 3572 -215 3576 -142
rect 3438 -228 3442 -224
rect 3473 -228 3477 -224
rect 3506 -228 3510 -224
rect 3539 -228 3543 -224
rect 3572 -228 3576 -224
rect 2235 -304 2239 -297
rect 2281 -304 2285 -297
rect 2326 -304 2330 -297
rect 2369 -304 2373 -297
rect 2414 -304 2418 -297
rect 2457 -304 2461 -297
rect 2617 -304 2621 -297
rect 2663 -304 2667 -297
rect 2708 -304 2712 -297
rect 2751 -304 2755 -297
rect 2796 -304 2800 -297
rect 2839 -304 2843 -297
rect 2999 -304 3003 -297
rect 3045 -304 3049 -297
rect 3090 -304 3094 -297
rect 3133 -304 3137 -297
rect 3178 -304 3182 -297
rect 3221 -304 3225 -297
rect 2050 -324 2054 -321
rect 2082 -324 2086 -321
rect 2116 -324 2120 -321
rect -318 -362 -314 -356
rect -286 -362 -282 -358
rect -252 -362 -248 -358
rect -172 -361 -168 -355
rect -140 -361 -136 -357
rect -106 -361 -102 -357
rect -42 -358 -38 -352
rect -10 -358 -6 -354
rect 24 -358 28 -354
rect 99 -359 103 -353
rect 131 -359 135 -355
rect 165 -359 169 -355
rect -318 -405 -314 -371
rect -317 -410 -314 -405
rect -318 -420 -314 -410
rect -286 -420 -282 -371
rect -252 -420 -248 -371
rect -172 -404 -168 -370
rect -171 -409 -168 -404
rect -172 -419 -168 -409
rect -140 -419 -136 -370
rect -106 -419 -102 -370
rect -42 -401 -38 -367
rect -41 -406 -38 -401
rect -42 -416 -38 -406
rect -10 -416 -6 -367
rect 24 -416 28 -367
rect 99 -402 103 -368
rect 100 -407 103 -402
rect 99 -417 103 -407
rect 131 -417 135 -368
rect 165 -417 169 -368
rect -42 -428 -38 -425
rect -10 -428 -6 -425
rect 24 -428 28 -425
rect 410 -422 414 -416
rect 442 -422 446 -418
rect 476 -422 480 -418
rect -318 -432 -314 -429
rect -286 -432 -282 -429
rect -252 -432 -248 -429
rect -172 -431 -168 -428
rect -140 -431 -136 -428
rect -106 -431 -102 -428
rect 99 -429 103 -426
rect 131 -429 135 -426
rect 165 -429 169 -426
rect 410 -465 414 -431
rect 411 -470 414 -465
rect 410 -480 414 -470
rect 442 -480 446 -431
rect 476 -480 480 -431
rect 2102 -484 2203 -481
rect 410 -492 414 -489
rect 442 -492 446 -489
rect 476 -492 480 -489
rect 2067 -510 2070 -501
rect 2102 -510 2105 -484
rect 2137 -510 2140 -501
rect 2169 -510 2172 -501
rect 2200 -510 2203 -484
rect 2233 -510 2236 -501
rect -261 -528 -257 -522
rect -229 -528 -225 -524
rect -195 -528 -191 -524
rect -261 -571 -257 -537
rect -260 -576 -257 -571
rect -261 -586 -257 -576
rect -229 -586 -225 -537
rect -195 -586 -191 -537
rect -85 -584 -81 -578
rect -53 -584 -49 -580
rect -19 -584 -15 -580
rect -261 -598 -257 -595
rect -229 -598 -225 -595
rect -195 -598 -191 -595
rect -85 -627 -81 -593
rect -84 -632 -81 -627
rect -85 -642 -81 -632
rect -53 -642 -49 -593
rect -19 -642 -15 -593
rect 169 -594 173 -588
rect 201 -594 205 -590
rect 235 -594 239 -590
rect 2067 -599 2070 -516
rect 2102 -599 2105 -516
rect 2137 -599 2140 -516
rect 2169 -599 2172 -516
rect 2200 -599 2203 -516
rect 2233 -599 2236 -516
rect 169 -637 173 -603
rect 170 -642 173 -637
rect -85 -654 -81 -651
rect -53 -654 -49 -651
rect -19 -654 -15 -651
rect 169 -652 173 -642
rect 201 -652 205 -603
rect 235 -652 239 -603
rect 2067 -616 2070 -605
rect 2102 -613 2105 -605
rect 2137 -616 2140 -605
rect 2169 -613 2172 -605
rect 2200 -613 2203 -605
rect 2233 -613 2236 -605
rect 2067 -618 2140 -616
rect 169 -664 173 -661
rect 201 -664 205 -661
rect 235 -664 239 -661
rect 2101 -731 2202 -728
rect 2066 -757 2069 -748
rect 2101 -757 2104 -731
rect 2136 -757 2139 -748
rect 2168 -757 2171 -748
rect 2199 -757 2202 -731
rect 2232 -757 2235 -748
rect 2066 -846 2069 -763
rect 2101 -846 2104 -763
rect 2136 -846 2139 -763
rect 2168 -846 2171 -763
rect 2199 -846 2202 -763
rect 2232 -846 2235 -763
rect 2426 -803 2430 -798
rect 2472 -803 2476 -798
rect 2517 -803 2521 -798
rect 2560 -803 2564 -798
rect 2605 -803 2609 -798
rect 2648 -803 2652 -798
rect 2066 -863 2069 -852
rect 2101 -860 2104 -852
rect 2136 -863 2139 -852
rect 2168 -860 2171 -852
rect 2199 -860 2202 -852
rect 2232 -860 2235 -852
rect 2066 -865 2139 -863
rect 2426 -906 2430 -814
rect 2472 -861 2476 -814
rect 2471 -870 2476 -861
rect 2517 -862 2521 -814
rect 2560 -862 2564 -814
rect 2472 -906 2476 -870
rect 2519 -871 2521 -862
rect 2562 -871 2564 -862
rect 2605 -864 2609 -814
rect 2517 -906 2521 -871
rect 2560 -906 2564 -871
rect 2606 -873 2609 -864
rect 2605 -906 2609 -873
rect 2648 -906 2652 -814
rect 2426 -924 2430 -917
rect 2472 -924 2476 -917
rect 2517 -924 2521 -917
rect 2560 -924 2564 -917
rect 2605 -924 2609 -917
rect 2648 -924 2652 -917
rect 2105 -957 2206 -954
rect 2070 -983 2073 -974
rect 2105 -983 2108 -957
rect 2140 -983 2143 -974
rect 2172 -983 2175 -974
rect 2203 -983 2206 -957
rect 2236 -983 2239 -974
rect 2070 -1072 2073 -989
rect 2105 -1072 2108 -989
rect 2140 -1072 2143 -989
rect 2172 -1072 2175 -989
rect 2203 -1072 2206 -989
rect 2236 -1072 2239 -989
rect 2070 -1089 2073 -1078
rect 2105 -1086 2108 -1078
rect 2140 -1089 2143 -1078
rect 2172 -1086 2175 -1078
rect 2203 -1086 2206 -1078
rect 2236 -1086 2239 -1078
rect 2070 -1091 2143 -1089
rect 2102 -1164 2203 -1161
rect 2067 -1190 2070 -1181
rect 2102 -1190 2105 -1164
rect 2137 -1190 2140 -1181
rect 2169 -1190 2172 -1181
rect 2200 -1190 2203 -1164
rect 2233 -1190 2236 -1181
rect 2067 -1279 2070 -1196
rect 2102 -1279 2105 -1196
rect 2137 -1279 2140 -1196
rect 2169 -1279 2172 -1196
rect 2200 -1279 2203 -1196
rect 2233 -1279 2236 -1196
rect 2067 -1296 2070 -1285
rect 2102 -1293 2105 -1285
rect 2137 -1296 2140 -1285
rect 2169 -1293 2172 -1285
rect 2200 -1293 2203 -1285
rect 2233 -1293 2236 -1285
rect 2067 -1298 2140 -1296
rect 2093 -1399 2097 -1393
rect 2125 -1399 2129 -1395
rect 2159 -1399 2163 -1395
rect 2093 -1442 2097 -1408
rect 2094 -1447 2097 -1442
rect 2093 -1457 2097 -1447
rect 2125 -1457 2129 -1408
rect 2159 -1457 2163 -1408
rect 2286 -1409 2290 -1404
rect 2332 -1409 2336 -1404
rect 2377 -1409 2381 -1404
rect 2420 -1409 2424 -1404
rect 2465 -1409 2469 -1404
rect 2508 -1409 2512 -1404
rect 2658 -1408 2662 -1403
rect 2704 -1408 2708 -1403
rect 2749 -1408 2753 -1403
rect 2792 -1408 2796 -1403
rect 2837 -1408 2841 -1403
rect 2880 -1408 2884 -1403
rect 3032 -1408 3036 -1403
rect 3078 -1408 3082 -1403
rect 3123 -1408 3127 -1403
rect 3166 -1408 3170 -1403
rect 3211 -1408 3215 -1403
rect 3254 -1408 3258 -1403
rect 2093 -1469 2097 -1466
rect 2125 -1469 2129 -1466
rect 2159 -1469 2163 -1466
rect 2286 -1512 2290 -1420
rect 2332 -1467 2336 -1420
rect 2331 -1476 2336 -1467
rect 2377 -1468 2381 -1420
rect 2420 -1468 2424 -1420
rect 2332 -1512 2336 -1476
rect 2379 -1477 2381 -1468
rect 2422 -1477 2424 -1468
rect 2465 -1470 2469 -1420
rect 2377 -1512 2381 -1477
rect 2420 -1512 2424 -1477
rect 2466 -1479 2469 -1470
rect 2465 -1512 2469 -1479
rect 2508 -1512 2512 -1420
rect 2658 -1511 2662 -1419
rect 2704 -1466 2708 -1419
rect 2703 -1475 2708 -1466
rect 2749 -1467 2753 -1419
rect 2792 -1467 2796 -1419
rect 2704 -1511 2708 -1475
rect 2751 -1476 2753 -1467
rect 2794 -1476 2796 -1467
rect 2837 -1469 2841 -1419
rect 2749 -1511 2753 -1476
rect 2792 -1511 2796 -1476
rect 2838 -1478 2841 -1469
rect 2837 -1511 2841 -1478
rect 2880 -1511 2884 -1419
rect 3032 -1511 3036 -1419
rect 3078 -1466 3082 -1419
rect 3077 -1475 3082 -1466
rect 3123 -1467 3127 -1419
rect 3166 -1467 3170 -1419
rect 3078 -1511 3082 -1475
rect 3125 -1476 3127 -1467
rect 3168 -1476 3170 -1467
rect 3211 -1469 3215 -1419
rect 3123 -1511 3127 -1476
rect 3166 -1511 3170 -1476
rect 3212 -1478 3215 -1469
rect 3211 -1511 3215 -1478
rect 3254 -1511 3258 -1419
rect 3488 -1460 3492 -1450
rect 3523 -1460 3527 -1450
rect 3556 -1460 3560 -1450
rect 3589 -1460 3593 -1450
rect 3622 -1460 3626 -1450
rect 2128 -1525 2132 -1513
rect 2286 -1530 2290 -1523
rect 2332 -1530 2336 -1523
rect 2377 -1530 2381 -1523
rect 2420 -1530 2424 -1523
rect 2465 -1530 2469 -1523
rect 2508 -1530 2512 -1523
rect 2658 -1529 2662 -1522
rect 2704 -1529 2708 -1522
rect 2749 -1529 2753 -1522
rect 2792 -1529 2796 -1522
rect 2837 -1529 2841 -1522
rect 2880 -1529 2884 -1522
rect 3032 -1529 3036 -1522
rect 3078 -1529 3082 -1522
rect 3123 -1529 3127 -1522
rect 3166 -1529 3170 -1522
rect 3211 -1529 3215 -1522
rect 3254 -1529 3258 -1522
rect 2128 -1563 2132 -1535
rect 3488 -1542 3492 -1469
rect 3523 -1542 3527 -1469
rect 3556 -1542 3560 -1469
rect 3589 -1542 3593 -1469
rect 3622 -1542 3626 -1469
rect 3488 -1555 3492 -1551
rect 3523 -1555 3527 -1551
rect 3556 -1555 3560 -1551
rect 3589 -1555 3593 -1551
rect 3622 -1555 3626 -1551
rect 2325 -1571 2329 -1559
rect 2128 -1592 2132 -1577
rect 2325 -1609 2329 -1581
rect 2733 -1595 2737 -1583
rect 3160 -1594 3164 -1582
rect 2325 -1638 2329 -1623
rect 2733 -1633 2737 -1605
rect 3160 -1632 3164 -1604
rect 2733 -1662 2737 -1647
rect 3160 -1661 3164 -1646
<< polycontact >>
rect 498 1998 503 2003
rect 527 1997 532 2002
rect 617 2007 621 2012
rect 646 1980 651 1986
rect 716 1998 721 2003
rect 745 1997 750 2002
rect 835 2007 839 2012
rect 864 1980 869 1986
rect 949 2000 954 2005
rect 978 1999 983 2004
rect 1068 2009 1072 2014
rect 1097 1982 1102 1988
rect 1209 2001 1214 2006
rect 1238 2000 1243 2005
rect 1328 2010 1332 2015
rect 1357 1983 1362 1989
rect 527 1800 532 1805
rect 556 1799 561 1804
rect 646 1809 650 1814
rect 675 1782 680 1788
rect 756 1795 760 1800
rect 787 1795 791 1800
rect 819 1808 825 1814
rect 1153 1797 1158 1802
rect 929 1787 933 1791
rect 947 1789 951 1793
rect 966 1790 970 1794
rect 1182 1796 1187 1801
rect 1272 1806 1276 1811
rect 1301 1779 1306 1785
rect 1382 1792 1386 1797
rect 1413 1792 1417 1797
rect 1445 1805 1451 1811
rect 1753 1797 1758 1802
rect 1555 1784 1559 1788
rect 1573 1786 1577 1790
rect 1592 1787 1596 1791
rect 1782 1796 1787 1801
rect 1872 1806 1876 1811
rect 1901 1779 1906 1785
rect 1982 1792 1986 1797
rect 2013 1792 2017 1797
rect 2045 1805 2051 1811
rect 2356 1800 2361 1805
rect 2155 1784 2159 1788
rect 2173 1786 2177 1790
rect 2192 1787 2196 1791
rect 2385 1799 2390 1804
rect 2475 1809 2479 1814
rect 2504 1782 2509 1788
rect 2585 1795 2589 1800
rect 2616 1795 2620 1800
rect 2648 1808 2654 1814
rect 2758 1787 2762 1791
rect 2776 1789 2780 1793
rect 2795 1790 2799 1794
rect 772 1656 776 1661
rect 803 1656 807 1661
rect 835 1669 841 1675
rect 1398 1653 1402 1658
rect 1429 1653 1433 1658
rect 1461 1666 1467 1672
rect 1998 1653 2002 1658
rect 2029 1653 2033 1658
rect 2061 1666 2067 1672
rect 2601 1656 2605 1661
rect 2632 1656 2636 1661
rect 2664 1669 2670 1675
rect 537 1544 542 1549
rect 566 1543 571 1548
rect 656 1553 660 1558
rect 685 1526 690 1532
rect 1163 1541 1168 1546
rect 1192 1540 1197 1545
rect 1282 1550 1286 1555
rect 1311 1523 1316 1529
rect 1763 1541 1768 1546
rect 1792 1540 1797 1545
rect 1882 1550 1886 1555
rect 1911 1523 1916 1529
rect 2366 1544 2371 1549
rect 2395 1543 2400 1548
rect 2485 1553 2489 1558
rect 2514 1526 2519 1532
rect 551 1183 556 1188
rect 580 1182 585 1187
rect 670 1192 674 1197
rect 699 1165 704 1171
rect 769 1183 774 1188
rect 798 1182 803 1187
rect 888 1192 892 1197
rect 917 1165 922 1171
rect 1002 1185 1007 1190
rect 1031 1184 1036 1189
rect 1121 1194 1125 1199
rect 1150 1167 1155 1173
rect 1262 1186 1267 1191
rect 1291 1185 1296 1190
rect 1381 1195 1385 1200
rect 1410 1168 1415 1174
rect -404 1028 -400 1033
rect -373 1028 -369 1033
rect -341 1041 -335 1047
rect -268 1029 -264 1034
rect -237 1029 -233 1034
rect -205 1042 -199 1048
rect -133 1030 -129 1035
rect -102 1030 -98 1035
rect -70 1043 -64 1049
rect 4 1028 8 1033
rect 35 1028 39 1033
rect 67 1041 73 1047
rect 580 985 585 990
rect -405 908 -401 913
rect -374 908 -370 913
rect -342 921 -336 927
rect -259 909 -255 914
rect -228 909 -224 914
rect -196 922 -190 928
rect -129 912 -125 917
rect -98 912 -94 917
rect -66 925 -60 931
rect 609 984 614 989
rect 699 994 703 999
rect 728 967 733 973
rect 809 980 813 985
rect 840 980 844 985
rect 872 993 878 999
rect 1206 982 1211 987
rect 982 972 986 976
rect 1000 974 1004 978
rect 1019 975 1023 979
rect 12 911 16 916
rect 43 911 47 916
rect 75 924 81 930
rect 1235 981 1240 986
rect 1325 991 1329 996
rect 1354 964 1359 970
rect 1435 977 1439 982
rect 1466 977 1470 982
rect 1498 990 1504 996
rect 1806 982 1811 987
rect 1608 969 1612 973
rect 1626 971 1630 975
rect 1645 972 1649 976
rect 1835 981 1840 986
rect 1925 991 1929 996
rect 1954 964 1959 970
rect 2035 977 2039 982
rect 2066 977 2070 982
rect 2098 990 2104 996
rect 2409 985 2414 990
rect 2208 969 2212 973
rect 2226 971 2230 975
rect 2245 972 2249 976
rect 2438 984 2443 989
rect 2528 994 2532 999
rect 2557 967 2562 973
rect 2638 980 2642 985
rect 2669 980 2673 985
rect 2701 993 2707 999
rect 2811 972 2815 976
rect 2829 974 2833 978
rect 2848 975 2852 979
rect 825 841 829 846
rect 856 841 860 846
rect 888 854 894 860
rect 1451 838 1455 843
rect 1482 838 1486 843
rect 1514 851 1520 857
rect 2051 838 2055 843
rect 2082 838 2086 843
rect 2114 851 2120 857
rect 2654 841 2658 846
rect 2685 841 2689 846
rect 2717 854 2723 860
rect 590 729 595 734
rect 619 728 624 733
rect 709 738 713 743
rect 738 711 743 717
rect 1216 726 1221 731
rect 1245 725 1250 730
rect 1335 735 1339 740
rect 1364 708 1369 714
rect 1816 726 1821 731
rect 1845 725 1850 730
rect 1935 735 1939 740
rect 1964 708 1969 714
rect 2419 729 2424 734
rect 2448 728 2453 733
rect 2538 738 2542 743
rect 2567 711 2572 717
rect -385 585 -381 590
rect -354 585 -350 590
rect -322 598 -316 604
rect -249 586 -245 591
rect -218 586 -214 591
rect -186 599 -180 605
rect -114 587 -110 592
rect -83 587 -79 592
rect -51 600 -45 606
rect 23 585 27 590
rect 54 585 58 590
rect 86 598 92 604
rect -386 465 -382 470
rect -355 465 -351 470
rect -323 478 -317 484
rect -240 466 -236 471
rect -209 466 -205 471
rect -177 479 -171 485
rect -110 469 -106 474
rect -79 469 -75 474
rect -47 482 -41 488
rect 31 468 35 473
rect 62 468 66 473
rect -1221 405 -1215 409
rect -1046 411 -1042 416
rect -1015 411 -1011 416
rect -983 424 -977 430
rect 94 481 100 487
rect -1044 310 -1040 315
rect -1013 310 -1009 315
rect -981 323 -975 329
rect -1041 211 -1037 216
rect -1010 211 -1006 216
rect -978 224 -972 230
rect -1223 186 -1217 190
rect -372 160 -368 165
rect -341 160 -337 165
rect -309 173 -303 179
rect -236 161 -232 166
rect -205 161 -201 166
rect -173 174 -167 180
rect -101 162 -97 167
rect -70 162 -66 167
rect -38 175 -32 181
rect 36 160 40 165
rect 67 160 71 165
rect -1039 103 -1035 108
rect -1008 103 -1004 108
rect -976 116 -970 122
rect 99 173 105 179
rect -373 40 -369 45
rect -342 40 -338 45
rect -310 53 -304 59
rect -227 41 -223 46
rect -196 41 -192 46
rect -164 54 -158 60
rect -97 44 -93 49
rect -66 44 -62 49
rect -34 57 -28 63
rect 44 43 48 48
rect 75 43 79 48
rect 107 56 113 62
rect 2095 -11 2101 -7
rect 2365 -16 2371 -12
rect 2620 -10 2626 -6
rect 2888 -10 2894 -6
rect 3434 -181 3438 -177
rect -320 -290 -316 -285
rect -289 -290 -285 -285
rect -257 -277 -251 -271
rect -184 -289 -180 -284
rect -153 -289 -149 -284
rect -121 -276 -115 -270
rect -49 -288 -45 -283
rect -18 -288 -14 -283
rect 14 -275 20 -269
rect 88 -290 92 -285
rect 119 -290 123 -285
rect 151 -277 157 -271
rect 2226 -249 2235 -240
rect 2047 -302 2051 -297
rect 2078 -302 2082 -297
rect 2110 -289 2116 -283
rect 2271 -250 2280 -241
rect 2319 -251 2328 -242
rect 2362 -251 2371 -242
rect 2406 -253 2415 -244
rect 2447 -245 2457 -236
rect 2608 -249 2617 -240
rect 2653 -250 2662 -241
rect 2701 -251 2710 -242
rect 2744 -251 2753 -242
rect 2788 -253 2797 -244
rect 2829 -245 2839 -236
rect 2990 -249 2999 -240
rect 3035 -250 3044 -241
rect 3083 -251 3092 -242
rect 3126 -251 3135 -242
rect 3170 -253 3179 -244
rect 3211 -245 3221 -236
rect 3469 -182 3473 -178
rect 3502 -183 3506 -179
rect 3535 -184 3539 -180
rect 3567 -182 3572 -178
rect -321 -410 -317 -405
rect -290 -410 -286 -405
rect -258 -397 -252 -391
rect -175 -409 -171 -404
rect -144 -409 -140 -404
rect -112 -396 -106 -390
rect -45 -406 -41 -401
rect -14 -406 -10 -401
rect 18 -393 24 -387
rect 96 -407 100 -402
rect 127 -407 131 -402
rect 159 -394 165 -388
rect 407 -470 411 -465
rect 438 -470 442 -465
rect 470 -457 476 -451
rect -264 -576 -260 -571
rect -233 -576 -229 -571
rect -201 -563 -195 -557
rect 2060 -554 2067 -548
rect -88 -632 -84 -627
rect -57 -632 -53 -627
rect -25 -619 -19 -613
rect 2096 -555 2102 -549
rect 2163 -555 2169 -549
rect 2227 -579 2233 -574
rect 166 -642 170 -637
rect 197 -642 201 -637
rect 229 -629 235 -623
rect 2059 -801 2066 -795
rect 2095 -802 2101 -796
rect 2162 -802 2168 -796
rect 2226 -826 2232 -821
rect 2417 -869 2426 -860
rect 2462 -870 2471 -861
rect 2510 -871 2519 -862
rect 2553 -871 2562 -862
rect 2597 -873 2606 -864
rect 2638 -865 2648 -856
rect 2063 -1027 2070 -1021
rect 2099 -1028 2105 -1022
rect 2166 -1028 2172 -1022
rect 2230 -1052 2236 -1047
rect 2060 -1234 2067 -1228
rect 2096 -1235 2102 -1229
rect 2163 -1235 2169 -1229
rect 2227 -1259 2233 -1254
rect 2090 -1447 2094 -1442
rect 2121 -1447 2125 -1442
rect 2153 -1434 2159 -1428
rect 2277 -1475 2286 -1466
rect 2322 -1476 2331 -1467
rect 2370 -1477 2379 -1468
rect 2413 -1477 2422 -1468
rect 2457 -1479 2466 -1470
rect 2498 -1471 2508 -1462
rect 2649 -1474 2658 -1465
rect 2694 -1475 2703 -1466
rect 2742 -1476 2751 -1467
rect 2785 -1476 2794 -1467
rect 2829 -1478 2838 -1469
rect 2870 -1470 2880 -1461
rect 3023 -1474 3032 -1465
rect 3068 -1475 3077 -1466
rect 3116 -1476 3125 -1467
rect 3159 -1476 3168 -1467
rect 3203 -1478 3212 -1469
rect 3244 -1470 3254 -1461
rect 3484 -1508 3488 -1504
rect 2122 -1550 2128 -1546
rect 3519 -1509 3523 -1505
rect 3552 -1510 3556 -1506
rect 3585 -1511 3589 -1507
rect 3617 -1509 3622 -1505
rect 2319 -1596 2325 -1592
rect 2727 -1620 2733 -1616
rect 3154 -1619 3160 -1615
<< metal1 >>
rect 1176 2069 1195 2070
rect 939 2068 1387 2069
rect 888 2067 1387 2068
rect 459 2063 1387 2067
rect 459 2062 1127 2063
rect 459 2061 963 2062
rect -711 2060 466 2061
rect 488 2060 894 2061
rect -1290 2049 466 2060
rect -1290 2048 -701 2049
rect -1290 1245 -1275 2048
rect 460 1868 466 2049
rect 494 2041 498 2060
rect 523 2041 527 2060
rect 552 2041 556 2060
rect 581 2041 585 2060
rect 602 2046 643 2050
rect 602 2041 606 2046
rect 610 2041 614 2046
rect 639 2041 643 2046
rect 712 2041 716 2060
rect 741 2041 745 2060
rect 770 2041 774 2060
rect 799 2041 803 2060
rect 820 2046 861 2050
rect 820 2041 824 2046
rect 828 2041 832 2046
rect 857 2041 861 2046
rect 945 2043 949 2061
rect 974 2043 978 2062
rect 1003 2043 1007 2062
rect 1032 2043 1036 2062
rect 1053 2048 1094 2052
rect 1053 2043 1057 2048
rect 1061 2043 1065 2048
rect 1090 2043 1094 2048
rect 1205 2044 1209 2063
rect 1234 2044 1238 2063
rect 1263 2044 1267 2063
rect 1292 2044 1296 2063
rect 1313 2049 1354 2053
rect 1313 2044 1317 2049
rect 1321 2044 1325 2049
rect 1350 2044 1354 2049
rect 495 1998 498 2003
rect 515 1969 519 2037
rect 522 1997 527 2002
rect 522 1988 525 1997
rect 544 1986 548 2037
rect 573 2030 577 2037
rect 602 2030 606 2037
rect 573 2027 606 2030
rect 631 2030 635 2037
rect 660 2030 664 2037
rect 631 2027 664 2030
rect 609 2008 617 2012
rect 614 2007 617 2008
rect 660 2004 664 2027
rect 660 2003 675 2004
rect 660 1994 666 2003
rect 715 1998 716 2003
rect 544 1981 646 1986
rect 544 1969 548 1981
rect 642 1980 646 1981
rect 660 1977 664 1994
rect 602 1969 606 1970
rect 660 1969 664 1972
rect 733 1969 737 2037
rect 740 1997 745 2002
rect 741 1985 744 1997
rect 762 1986 766 2037
rect 791 2030 795 2037
rect 820 2030 824 2037
rect 791 2027 824 2030
rect 849 2030 853 2037
rect 878 2030 882 2037
rect 849 2027 882 2030
rect 827 2008 835 2012
rect 832 2007 835 2008
rect 762 1981 864 1986
rect 762 1969 766 1981
rect 860 1980 864 1981
rect 878 1977 882 2027
rect 946 2000 949 2005
rect 820 1969 824 1970
rect 878 1969 882 1972
rect 966 1971 970 2039
rect 973 1999 978 2004
rect 975 1987 978 1999
rect 995 1988 999 2039
rect 1024 2032 1028 2039
rect 1053 2032 1057 2039
rect 1024 2029 1057 2032
rect 1082 2032 1086 2039
rect 1111 2032 1115 2039
rect 1082 2029 1115 2032
rect 1060 2010 1068 2014
rect 1065 2009 1068 2010
rect 1111 2006 1115 2029
rect 1111 1996 1147 2006
rect 1206 2001 1209 2006
rect 995 1983 1097 1988
rect 995 1971 999 1983
rect 1093 1982 1097 1983
rect 1111 1979 1115 1996
rect 1053 1971 1057 1972
rect 1111 1971 1115 1974
rect 1226 1972 1230 2040
rect 1233 2000 1238 2005
rect 1234 1989 1237 2000
rect 1255 1989 1259 2040
rect 1284 2033 1288 2040
rect 1313 2033 1317 2040
rect 1284 2030 1317 2033
rect 1342 2033 1346 2040
rect 1371 2033 1375 2040
rect 1342 2030 1375 2033
rect 1320 2011 1328 2015
rect 1325 2010 1328 2011
rect 1371 2007 1375 2030
rect 1371 2006 1379 2007
rect 1371 1998 1420 2006
rect 1371 1997 1379 1998
rect 1255 1984 1357 1989
rect 1255 1972 1259 1984
rect 1353 1983 1357 1984
rect 1371 1980 1375 1997
rect 1313 1972 1317 1973
rect 1371 1972 1375 1975
rect 577 1965 581 1969
rect 635 1965 639 1969
rect 795 1965 799 1969
rect 853 1965 857 1969
rect 1028 1967 1032 1971
rect 1086 1967 1090 1971
rect 1288 1968 1292 1972
rect 1346 1968 1350 1972
rect 494 1961 498 1965
rect 523 1961 527 1965
rect 552 1961 556 1965
rect 610 1961 614 1965
rect 712 1961 716 1965
rect 741 1961 745 1965
rect 770 1961 774 1965
rect 828 1961 832 1965
rect 945 1963 949 1967
rect 974 1963 978 1967
rect 1003 1963 1007 1967
rect 1061 1963 1065 1967
rect 942 1962 1130 1963
rect 891 1961 1200 1962
rect 1205 1961 1209 1968
rect 1234 1964 1238 1968
rect 1263 1964 1267 1968
rect 1321 1964 1325 1968
rect 1212 1963 1390 1964
rect 1212 1961 2937 1963
rect 495 1957 2937 1961
rect 495 1956 1221 1957
rect 1382 1956 2937 1957
rect 495 1955 946 1956
rect 495 1954 897 1955
rect 460 1862 730 1868
rect 1187 1865 1191 1866
rect 1086 1862 1356 1865
rect 460 1861 533 1862
rect -303 1805 -293 1806
rect -303 1801 443 1805
rect -303 1765 -293 1801
rect 460 1620 474 1861
rect 523 1843 527 1861
rect 552 1843 556 1862
rect 581 1843 585 1862
rect 610 1843 614 1862
rect 725 1859 730 1862
rect 975 1859 1356 1862
rect 725 1858 1159 1859
rect 725 1853 1100 1858
rect 725 1852 998 1853
rect 631 1848 672 1852
rect 631 1843 635 1848
rect 639 1843 643 1848
rect 668 1843 672 1848
rect 750 1843 755 1852
rect 781 1843 786 1852
rect 814 1843 819 1852
rect 544 1815 548 1839
rect 544 1811 564 1815
rect 525 1800 527 1805
rect 544 1771 548 1811
rect 573 1788 577 1839
rect 602 1832 606 1839
rect 631 1832 635 1839
rect 602 1829 635 1832
rect 660 1832 664 1839
rect 689 1832 693 1839
rect 660 1829 693 1832
rect 638 1810 646 1814
rect 643 1809 646 1810
rect 689 1806 693 1829
rect 769 1814 774 1838
rect 800 1814 805 1838
rect 769 1808 819 1814
rect 689 1803 697 1806
rect 689 1798 731 1803
rect 689 1796 697 1798
rect 573 1783 675 1788
rect 573 1771 577 1783
rect 671 1782 675 1783
rect 689 1779 693 1796
rect 631 1771 635 1772
rect 689 1771 693 1774
rect 606 1767 610 1771
rect 664 1767 668 1771
rect 523 1763 527 1767
rect 552 1763 556 1767
rect 581 1764 585 1767
rect 579 1763 585 1764
rect 639 1763 643 1767
rect 495 1756 701 1763
rect 495 1507 507 1756
rect 724 1661 731 1798
rect 755 1795 756 1800
rect 786 1795 787 1800
rect 800 1785 805 1808
rect 833 1785 838 1838
rect 992 1829 998 1852
rect 912 1824 998 1829
rect 926 1818 930 1824
rect 963 1818 967 1824
rect 940 1814 944 1818
rect 954 1794 958 1814
rect 973 1800 977 1814
rect 774 1780 781 1785
rect 907 1787 929 1791
rect 946 1789 947 1793
rect 954 1790 966 1794
rect 973 1793 976 1800
rect 907 1786 928 1787
rect 750 1776 755 1780
rect 814 1776 819 1780
rect 744 1775 845 1776
rect 751 1769 845 1775
rect 759 1713 888 1720
rect 766 1704 771 1713
rect 797 1704 802 1713
rect 830 1704 835 1713
rect 785 1675 790 1699
rect 816 1675 821 1699
rect 785 1669 835 1675
rect 849 1672 854 1699
rect 907 1672 914 1786
rect 954 1785 958 1790
rect 936 1782 958 1785
rect 936 1777 940 1782
rect 954 1777 958 1782
rect 973 1777 977 1793
rect 926 1770 930 1773
rect 944 1770 948 1773
rect 963 1770 967 1773
rect 922 1769 986 1770
rect 931 1767 986 1769
rect 991 1720 998 1824
rect 954 1713 998 1720
rect 724 1656 772 1661
rect 800 1656 803 1661
rect 535 1607 715 1613
rect 527 1606 715 1607
rect 533 1587 537 1606
rect 562 1587 566 1606
rect 591 1587 595 1606
rect 620 1587 624 1606
rect 641 1592 682 1596
rect 641 1587 645 1592
rect 649 1587 653 1592
rect 678 1587 682 1592
rect 534 1544 537 1549
rect 554 1515 558 1583
rect 583 1532 587 1583
rect 612 1576 616 1583
rect 641 1576 645 1583
rect 612 1573 645 1576
rect 670 1576 674 1583
rect 699 1576 703 1583
rect 670 1573 703 1576
rect 648 1554 656 1558
rect 653 1553 656 1554
rect 699 1550 703 1573
rect 699 1540 707 1550
rect 583 1527 685 1532
rect 583 1515 587 1527
rect 681 1526 685 1527
rect 699 1523 703 1540
rect 641 1515 645 1516
rect 699 1515 703 1518
rect 616 1511 620 1515
rect 674 1511 678 1515
rect 533 1507 537 1511
rect 562 1507 566 1511
rect 591 1507 595 1511
rect 649 1507 653 1511
rect 495 1500 718 1507
rect 495 1450 507 1500
rect 724 1479 731 1656
rect 816 1646 821 1669
rect 849 1667 914 1672
rect 849 1646 854 1667
rect 790 1641 797 1646
rect 766 1637 771 1641
rect 830 1637 835 1641
rect 568 1472 731 1479
rect 760 1630 867 1637
rect 158 1442 507 1450
rect 760 1442 774 1630
rect 1086 1617 1100 1853
rect 1149 1840 1153 1858
rect 1178 1840 1182 1859
rect 1207 1840 1211 1859
rect 1236 1840 1240 1859
rect 1351 1856 1356 1859
rect 1686 1859 1956 1865
rect 1686 1858 1759 1859
rect 1686 1857 1700 1858
rect 1619 1856 1700 1857
rect 1351 1849 1700 1856
rect 1257 1845 1298 1849
rect 1257 1840 1261 1845
rect 1265 1840 1269 1845
rect 1294 1840 1298 1845
rect 1376 1840 1381 1849
rect 1407 1840 1412 1849
rect 1440 1840 1445 1849
rect 1170 1812 1174 1836
rect 1170 1808 1190 1812
rect 1151 1797 1153 1802
rect 1170 1768 1174 1808
rect 1199 1785 1203 1836
rect 1228 1829 1232 1836
rect 1257 1829 1261 1836
rect 1228 1826 1261 1829
rect 1286 1829 1290 1836
rect 1315 1829 1319 1836
rect 1286 1826 1319 1829
rect 1264 1807 1272 1811
rect 1269 1806 1272 1807
rect 1315 1803 1319 1826
rect 1395 1811 1400 1835
rect 1426 1811 1431 1835
rect 1395 1805 1445 1811
rect 1315 1800 1323 1803
rect 1315 1795 1357 1800
rect 1315 1793 1323 1795
rect 1199 1780 1301 1785
rect 1199 1768 1203 1780
rect 1297 1779 1301 1780
rect 1315 1776 1319 1793
rect 1257 1768 1261 1769
rect 1315 1768 1319 1771
rect 1232 1764 1236 1768
rect 1290 1764 1294 1768
rect 1149 1760 1153 1764
rect 1178 1760 1182 1764
rect 1207 1760 1211 1764
rect 1265 1760 1269 1764
rect 1121 1753 1327 1760
rect 158 1439 774 1442
rect 1121 1504 1133 1753
rect 1350 1658 1357 1795
rect 1381 1792 1382 1797
rect 1412 1792 1413 1797
rect 1426 1782 1431 1805
rect 1459 1782 1464 1835
rect 1618 1826 1624 1849
rect 1538 1821 1624 1826
rect 1552 1815 1556 1821
rect 1589 1815 1593 1821
rect 1566 1811 1570 1815
rect 1580 1791 1584 1811
rect 1599 1794 1603 1811
rect 1400 1777 1407 1782
rect 1533 1784 1555 1788
rect 1572 1786 1573 1790
rect 1580 1787 1592 1791
rect 1599 1790 1606 1794
rect 1533 1783 1554 1784
rect 1376 1773 1381 1777
rect 1440 1773 1445 1777
rect 1370 1772 1471 1773
rect 1377 1766 1471 1772
rect 1385 1710 1514 1717
rect 1392 1701 1397 1710
rect 1423 1701 1428 1710
rect 1456 1701 1461 1710
rect 1411 1672 1416 1696
rect 1442 1672 1447 1696
rect 1411 1666 1461 1672
rect 1475 1669 1480 1696
rect 1533 1669 1540 1783
rect 1580 1782 1584 1787
rect 1562 1779 1584 1782
rect 1562 1774 1566 1779
rect 1580 1774 1584 1779
rect 1599 1774 1603 1790
rect 1552 1767 1556 1770
rect 1570 1767 1574 1770
rect 1589 1767 1593 1770
rect 1548 1766 1612 1767
rect 1557 1764 1612 1766
rect 1617 1717 1624 1821
rect 1580 1710 1624 1717
rect 1350 1653 1398 1658
rect 1426 1653 1429 1658
rect 1161 1604 1341 1610
rect 1153 1603 1341 1604
rect 1159 1584 1163 1603
rect 1188 1584 1192 1603
rect 1217 1584 1221 1603
rect 1246 1584 1250 1603
rect 1267 1589 1308 1593
rect 1267 1584 1271 1589
rect 1275 1584 1279 1589
rect 1304 1584 1308 1589
rect 1160 1541 1163 1546
rect 1180 1512 1184 1580
rect 1209 1529 1213 1580
rect 1238 1573 1242 1580
rect 1267 1573 1271 1580
rect 1238 1570 1271 1573
rect 1296 1573 1300 1580
rect 1325 1573 1329 1580
rect 1296 1570 1329 1573
rect 1274 1551 1282 1555
rect 1279 1550 1282 1551
rect 1325 1547 1329 1570
rect 1325 1537 1333 1547
rect 1209 1524 1311 1529
rect 1209 1512 1213 1524
rect 1307 1523 1311 1524
rect 1325 1520 1329 1537
rect 1267 1512 1271 1513
rect 1325 1512 1329 1515
rect 1242 1508 1246 1512
rect 1300 1508 1304 1512
rect 1159 1504 1163 1508
rect 1188 1504 1192 1508
rect 1217 1504 1221 1508
rect 1275 1504 1279 1508
rect 1121 1497 1344 1504
rect 1121 1439 1133 1497
rect 1350 1476 1357 1653
rect 1442 1643 1447 1666
rect 1475 1664 1540 1669
rect 1475 1643 1480 1664
rect 1416 1638 1423 1643
rect 1392 1634 1397 1638
rect 1456 1634 1461 1638
rect 1194 1469 1357 1476
rect 1386 1627 1493 1634
rect 1386 1439 1400 1627
rect 1686 1617 1700 1849
rect 1749 1840 1753 1858
rect 1778 1840 1782 1859
rect 1786 1858 1790 1859
rect 1807 1840 1811 1859
rect 1836 1840 1840 1859
rect 1951 1856 1956 1859
rect 2289 1862 2559 1868
rect 2289 1861 2362 1862
rect 1951 1851 2224 1856
rect 2289 1851 2303 1861
rect 1951 1849 2303 1851
rect 1857 1845 1898 1849
rect 1857 1840 1861 1845
rect 1865 1840 1869 1845
rect 1894 1840 1898 1845
rect 1976 1840 1981 1849
rect 2007 1840 2012 1849
rect 2040 1840 2045 1849
rect 2218 1843 2303 1849
rect 1770 1812 1774 1836
rect 1770 1808 1790 1812
rect 1751 1797 1753 1802
rect 1770 1768 1774 1808
rect 1799 1785 1803 1836
rect 1828 1829 1832 1836
rect 1857 1829 1861 1836
rect 1828 1826 1861 1829
rect 1886 1829 1890 1836
rect 1915 1829 1919 1836
rect 1886 1826 1919 1829
rect 1864 1807 1872 1811
rect 1869 1806 1872 1807
rect 1915 1803 1919 1826
rect 1995 1811 2000 1835
rect 2026 1811 2031 1835
rect 1995 1805 2045 1811
rect 1915 1800 1923 1803
rect 1915 1795 1957 1800
rect 1915 1793 1923 1795
rect 1799 1780 1901 1785
rect 1799 1768 1803 1780
rect 1897 1779 1901 1780
rect 1915 1776 1919 1793
rect 1857 1768 1861 1769
rect 1915 1768 1919 1771
rect 1832 1764 1836 1768
rect 1890 1764 1894 1768
rect 1749 1760 1753 1764
rect 1778 1760 1782 1764
rect 1807 1760 1811 1764
rect 1865 1760 1869 1764
rect 1721 1753 1927 1760
rect 158 1435 1400 1439
rect 1721 1504 1733 1753
rect 1950 1658 1957 1795
rect 1981 1792 1982 1797
rect 2012 1792 2013 1797
rect 2026 1782 2031 1805
rect 2059 1782 2064 1835
rect 2218 1826 2224 1843
rect 2138 1821 2224 1826
rect 2152 1815 2156 1821
rect 2189 1815 2193 1821
rect 2166 1811 2170 1815
rect 2180 1791 2184 1811
rect 2199 1794 2203 1811
rect 2000 1777 2007 1782
rect 2133 1784 2155 1788
rect 2172 1786 2173 1790
rect 2180 1787 2192 1791
rect 2199 1790 2206 1794
rect 2133 1783 2154 1784
rect 1976 1773 1981 1777
rect 2040 1773 2045 1777
rect 1970 1772 2071 1773
rect 1977 1766 2071 1772
rect 1985 1710 2114 1717
rect 1992 1701 1997 1710
rect 2023 1701 2028 1710
rect 2056 1701 2061 1710
rect 2011 1672 2016 1696
rect 2042 1672 2047 1696
rect 2011 1666 2061 1672
rect 2075 1669 2080 1696
rect 2133 1669 2140 1783
rect 2180 1782 2184 1787
rect 2162 1779 2184 1782
rect 2162 1774 2166 1779
rect 2180 1774 2184 1779
rect 2199 1774 2203 1790
rect 2152 1767 2156 1770
rect 2170 1767 2174 1770
rect 2189 1767 2193 1770
rect 2148 1766 2212 1767
rect 2157 1764 2212 1766
rect 2217 1717 2224 1821
rect 2180 1710 2224 1717
rect 1950 1653 1998 1658
rect 2026 1653 2029 1658
rect 1761 1604 1941 1610
rect 1753 1603 1941 1604
rect 1759 1584 1763 1603
rect 1788 1584 1792 1603
rect 1817 1584 1821 1603
rect 1846 1584 1850 1603
rect 1867 1589 1908 1593
rect 1867 1584 1871 1589
rect 1875 1584 1879 1589
rect 1904 1584 1908 1589
rect 1761 1541 1763 1546
rect 1780 1512 1784 1580
rect 1809 1529 1813 1580
rect 1838 1573 1842 1580
rect 1867 1573 1871 1580
rect 1838 1570 1871 1573
rect 1896 1573 1900 1580
rect 1925 1573 1929 1580
rect 1896 1570 1929 1573
rect 1874 1551 1882 1555
rect 1879 1550 1882 1551
rect 1925 1547 1929 1570
rect 1925 1537 1933 1547
rect 1809 1524 1911 1529
rect 1809 1512 1813 1524
rect 1907 1523 1911 1524
rect 1925 1520 1929 1537
rect 1867 1512 1871 1513
rect 1925 1512 1929 1515
rect 1842 1508 1846 1512
rect 1900 1508 1904 1512
rect 1759 1504 1763 1508
rect 1788 1504 1792 1508
rect 1817 1504 1821 1508
rect 1875 1504 1879 1508
rect 1721 1497 1944 1504
rect 1721 1439 1733 1497
rect 1950 1476 1957 1653
rect 2042 1643 2047 1666
rect 2075 1664 2140 1669
rect 2075 1643 2080 1664
rect 2016 1638 2023 1643
rect 1992 1634 1997 1638
rect 2056 1634 2061 1638
rect 1794 1469 1957 1476
rect 1986 1627 2093 1634
rect 1986 1439 2000 1627
rect 2289 1620 2303 1843
rect 2352 1843 2356 1861
rect 2381 1843 2385 1862
rect 2410 1843 2414 1862
rect 2439 1843 2443 1862
rect 2554 1859 2559 1862
rect 2554 1852 2827 1859
rect 2460 1848 2501 1852
rect 2460 1843 2464 1848
rect 2468 1843 2472 1848
rect 2497 1843 2501 1848
rect 2579 1843 2584 1852
rect 2610 1843 2615 1852
rect 2643 1843 2648 1852
rect 2373 1815 2377 1839
rect 2373 1811 2393 1815
rect 2354 1800 2356 1805
rect 2373 1771 2377 1811
rect 2402 1788 2406 1839
rect 2431 1832 2435 1839
rect 2460 1832 2464 1839
rect 2431 1829 2464 1832
rect 2489 1832 2493 1839
rect 2518 1832 2522 1839
rect 2489 1829 2522 1832
rect 2467 1810 2475 1814
rect 2472 1809 2475 1810
rect 2518 1806 2522 1829
rect 2598 1814 2603 1838
rect 2629 1814 2634 1838
rect 2598 1808 2648 1814
rect 2518 1803 2526 1806
rect 2518 1798 2560 1803
rect 2518 1796 2526 1798
rect 2402 1783 2504 1788
rect 2402 1771 2406 1783
rect 2500 1782 2504 1783
rect 2518 1779 2522 1796
rect 2460 1771 2464 1772
rect 2518 1771 2522 1774
rect 2435 1767 2439 1771
rect 2493 1767 2497 1771
rect 2352 1763 2356 1767
rect 2381 1763 2385 1767
rect 2410 1765 2414 1767
rect 2409 1763 2414 1765
rect 2468 1763 2472 1767
rect 2324 1756 2530 1763
rect 1721 1438 2000 1439
rect 2324 1507 2336 1756
rect 2553 1661 2560 1798
rect 2584 1795 2585 1800
rect 2615 1795 2616 1800
rect 2629 1785 2634 1808
rect 2662 1785 2667 1838
rect 2821 1829 2827 1852
rect 2741 1824 2827 1829
rect 2755 1818 2759 1824
rect 2792 1818 2796 1824
rect 2769 1814 2773 1818
rect 2783 1794 2787 1814
rect 2802 1797 2806 1814
rect 2603 1780 2610 1785
rect 2736 1787 2758 1791
rect 2775 1789 2776 1793
rect 2783 1790 2795 1794
rect 2802 1793 2811 1797
rect 2736 1786 2757 1787
rect 2579 1776 2584 1780
rect 2643 1776 2648 1780
rect 2573 1775 2674 1776
rect 2580 1769 2674 1775
rect 2588 1713 2717 1720
rect 2595 1704 2600 1713
rect 2626 1704 2631 1713
rect 2659 1704 2664 1713
rect 2614 1675 2619 1699
rect 2645 1675 2650 1699
rect 2614 1669 2664 1675
rect 2678 1672 2683 1699
rect 2736 1672 2743 1786
rect 2783 1785 2787 1790
rect 2765 1782 2787 1785
rect 2765 1777 2769 1782
rect 2783 1777 2787 1782
rect 2802 1777 2806 1793
rect 2755 1770 2759 1773
rect 2773 1770 2777 1773
rect 2792 1770 2796 1773
rect 2751 1769 2815 1770
rect 2760 1767 2815 1769
rect 2820 1720 2827 1824
rect 2783 1713 2827 1720
rect 2553 1656 2601 1661
rect 2629 1656 2632 1661
rect 2364 1607 2544 1613
rect 2356 1606 2544 1607
rect 2362 1587 2366 1606
rect 2391 1587 2395 1606
rect 2420 1587 2424 1606
rect 2449 1587 2453 1606
rect 2470 1592 2511 1596
rect 2470 1587 2474 1592
rect 2478 1587 2482 1592
rect 2507 1587 2511 1592
rect 2363 1544 2366 1549
rect 2383 1515 2387 1583
rect 2412 1532 2416 1583
rect 2441 1576 2445 1583
rect 2470 1576 2474 1583
rect 2441 1573 2474 1576
rect 2499 1576 2503 1583
rect 2528 1576 2532 1583
rect 2499 1573 2532 1576
rect 2477 1554 2485 1558
rect 2482 1553 2485 1554
rect 2528 1550 2532 1573
rect 2528 1540 2536 1550
rect 2412 1527 2514 1532
rect 2412 1515 2416 1527
rect 2510 1526 2514 1527
rect 2528 1523 2532 1540
rect 2470 1515 2474 1516
rect 2528 1515 2532 1518
rect 2445 1511 2449 1515
rect 2503 1511 2507 1515
rect 2362 1507 2366 1511
rect 2391 1507 2395 1511
rect 2420 1507 2424 1511
rect 2478 1507 2482 1511
rect 2324 1500 2547 1507
rect 2324 1442 2336 1500
rect 2553 1479 2560 1656
rect 2645 1646 2650 1669
rect 2678 1667 2743 1672
rect 2678 1646 2683 1667
rect 2619 1641 2626 1646
rect 2595 1637 2600 1641
rect 2659 1637 2664 1641
rect 2397 1472 2560 1479
rect 2589 1630 2696 1637
rect 2589 1442 2603 1630
rect 2324 1440 2603 1442
rect 2918 1440 2936 1956
rect 2324 1438 2936 1440
rect 1721 1435 2936 1438
rect 158 1434 2936 1435
rect 158 1421 171 1434
rect 506 1433 774 1434
rect 1121 1433 2936 1434
rect 1121 1430 2000 1433
rect 2577 1432 2936 1433
rect 159 1417 171 1421
rect 159 1374 172 1417
rect 992 1253 1440 1254
rect 941 1252 1440 1253
rect 512 1248 1440 1252
rect 512 1247 1180 1248
rect 512 1246 1016 1247
rect 512 1245 519 1246
rect 541 1245 947 1246
rect -1290 1244 -645 1245
rect -508 1244 519 1245
rect -1290 1235 519 1244
rect -1290 1096 -1275 1235
rect 475 1204 481 1235
rect -301 1102 -296 1140
rect -1291 1093 -437 1096
rect -1291 1092 -178 1093
rect -146 1092 -43 1094
rect -1291 1088 94 1092
rect -1291 1086 -1275 1088
rect -1291 816 -1281 1086
rect -1291 452 -1282 816
rect -778 651 -770 1088
rect -442 1087 94 1088
rect -442 1086 -178 1087
rect -652 1057 -470 1064
rect -459 1057 -458 1064
rect -542 1017 -519 1018
rect -537 1008 -519 1017
rect -537 1007 -501 1008
rect -442 972 -437 1086
rect -417 1085 -314 1086
rect -410 1076 -405 1085
rect -379 1076 -374 1085
rect -346 1076 -341 1085
rect -274 1077 -269 1086
rect -243 1077 -238 1086
rect -210 1077 -205 1086
rect -391 1047 -386 1071
rect -360 1047 -355 1071
rect -391 1041 -341 1047
rect -327 1045 -322 1071
rect -255 1048 -250 1072
rect -224 1048 -219 1072
rect -410 1028 -404 1033
rect -377 1028 -373 1033
rect -360 1018 -355 1041
rect -327 1039 -301 1045
rect -255 1042 -205 1048
rect -191 1046 -186 1072
rect -171 1046 -166 1075
rect -139 1078 -134 1087
rect -108 1078 -103 1087
rect -75 1078 -70 1087
rect -23 1086 94 1087
rect -9 1085 94 1086
rect -327 1018 -322 1039
rect -296 1029 -268 1034
rect -239 1029 -237 1034
rect -224 1019 -219 1042
rect -191 1040 -166 1046
rect -120 1049 -115 1073
rect -89 1049 -84 1073
rect -120 1043 -70 1049
rect -56 1047 -51 1073
rect -34 1047 -29 1078
rect -2 1076 3 1085
rect 29 1076 34 1085
rect 62 1076 67 1085
rect -191 1019 -186 1040
rect -136 1030 -133 1035
rect -104 1030 -102 1035
rect -89 1020 -84 1043
rect -56 1041 -29 1047
rect 17 1047 22 1071
rect 48 1047 53 1071
rect 17 1041 67 1047
rect -56 1020 -51 1041
rect 1 1028 4 1033
rect 33 1028 35 1033
rect -386 1013 -379 1018
rect -250 1014 -243 1019
rect -115 1015 -108 1020
rect 48 1018 53 1041
rect 81 1018 86 1071
rect -410 1009 -405 1013
rect -346 1009 -341 1013
rect -274 1010 -269 1014
rect -210 1010 -205 1014
rect -139 1011 -134 1015
rect -75 1011 -70 1015
rect 22 1013 29 1018
rect -280 1009 -167 1010
rect -145 1009 -32 1011
rect -2 1009 3 1013
rect 62 1009 67 1013
rect -416 1008 -303 1009
rect -280 1008 130 1009
rect -416 1007 130 1008
rect -417 1004 130 1007
rect -416 1003 -160 1004
rect -416 1002 -303 1003
rect -8 1002 130 1004
rect -142 975 -39 976
rect -173 973 102 975
rect -442 970 -315 972
rect -272 970 102 973
rect -442 969 102 970
rect -442 967 -169 969
rect -442 965 -315 967
rect -272 966 -169 967
rect -411 956 -406 965
rect -380 956 -375 965
rect -347 956 -342 965
rect -265 957 -260 966
rect -234 957 -229 966
rect -201 957 -196 966
rect -135 960 -130 969
rect -104 960 -99 969
rect -71 960 -66 969
rect -1 968 102 969
rect -392 927 -387 951
rect -361 927 -356 951
rect -392 921 -342 927
rect -328 925 -323 951
rect -246 928 -241 952
rect -215 928 -210 952
rect -409 908 -405 913
rect -376 908 -374 913
rect -361 898 -356 921
rect -328 919 -313 925
rect -246 922 -196 928
rect -182 925 -177 952
rect -116 931 -111 955
rect -85 931 -80 955
rect -116 925 -66 931
rect -52 929 -47 955
rect 6 959 11 968
rect 37 959 42 968
rect 70 959 75 968
rect 25 930 30 954
rect 56 930 61 954
rect -52 927 -43 929
rect -328 898 -323 919
rect -264 909 -259 914
rect -231 909 -228 914
rect -215 899 -210 922
rect -182 920 -170 925
rect -182 919 -163 920
rect -182 899 -177 919
rect -136 912 -129 917
rect -102 912 -98 917
rect -85 902 -80 925
rect -52 923 -36 927
rect -52 902 -47 923
rect 25 924 75 930
rect 89 929 94 954
rect 122 935 130 1002
rect 162 935 171 1191
rect 122 931 171 935
rect 89 928 107 929
rect -36 921 -31 922
rect 9 911 12 916
rect 39 911 43 916
rect -387 893 -380 898
rect -241 894 -234 899
rect -111 897 -104 902
rect 56 901 61 924
rect 89 923 102 928
rect 89 922 97 923
rect 89 901 94 922
rect -411 889 -406 893
rect -347 889 -342 893
rect -265 890 -260 894
rect -201 890 -196 894
rect -135 893 -130 897
rect -71 893 -66 897
rect 30 896 37 901
rect -141 891 -41 893
rect 6 892 11 896
rect 70 892 75 896
rect 122 892 130 931
rect -157 890 -41 891
rect 0 890 130 892
rect -317 889 130 890
rect -617 888 -590 889
rect -519 888 130 889
rect -617 886 130 888
rect -617 884 -137 886
rect 0 885 130 886
rect -617 882 -616 884
rect -602 883 -137 884
rect -602 882 -270 883
rect -135 874 -117 878
rect -122 659 -117 874
rect -779 650 -418 651
rect -779 649 -159 650
rect -127 649 -24 651
rect -779 644 113 649
rect -779 643 -159 644
rect -779 640 -418 643
rect -398 642 -295 643
rect -1096 468 -921 474
rect -1096 452 -1087 468
rect -1052 459 -1047 468
rect -1021 459 -1016 468
rect -988 459 -983 468
rect -1311 442 -1087 452
rect -1311 440 -1246 442
rect -1311 234 -1304 440
rect -1291 439 -1282 440
rect -1239 430 -1235 442
rect -1033 430 -1028 454
rect -1002 430 -997 454
rect -969 432 -964 454
rect -1191 411 -1187 426
rect -1033 424 -983 430
rect -1101 411 -1046 416
rect -1024 411 -1015 416
rect -1274 405 -1221 409
rect -1191 407 -1096 411
rect -1024 410 -1011 411
rect -1024 408 -1020 410
rect -1274 302 -1271 405
rect -1191 392 -1187 407
rect -1239 363 -1235 388
rect -1258 355 -1171 363
rect -1161 355 -1160 363
rect -1258 353 -1160 355
rect -1149 302 -1144 320
rect -1274 299 -1144 302
rect -1311 233 -1249 234
rect -1311 223 -1161 233
rect -1140 232 -1137 407
rect -1081 404 -1020 408
rect -1081 370 -1076 404
rect -1002 401 -997 424
rect -969 401 -964 424
rect -1028 396 -1021 401
rect -1052 392 -1047 396
rect -988 392 -983 396
rect -1058 385 -961 392
rect -929 373 -921 468
rect -778 433 -770 640
rect -1116 365 -1076 370
rect -1057 367 -921 373
rect -1116 315 -1111 365
rect -1050 358 -1045 367
rect -1019 358 -1014 367
rect -986 358 -981 367
rect -1031 329 -1026 353
rect -1000 329 -995 353
rect -1031 323 -981 329
rect -967 326 -962 353
rect -1116 310 -1044 315
rect -1241 211 -1237 223
rect -1278 186 -1223 190
rect -1193 189 -1189 207
rect -1116 189 -1111 310
rect -1017 310 -1013 315
rect -1017 309 -1009 310
rect -1000 300 -995 323
rect -967 300 -962 321
rect -1026 295 -1019 300
rect -1050 291 -1045 295
rect -986 291 -981 295
rect -1056 284 -958 291
rect -929 274 -921 367
rect -779 402 -770 433
rect -543 565 -511 575
rect -779 359 -771 402
rect -543 326 -540 565
rect -423 529 -418 640
rect -391 633 -386 642
rect -360 633 -355 642
rect -327 633 -322 642
rect -372 604 -367 628
rect -341 604 -336 628
rect -372 598 -322 604
rect -308 602 -303 628
rect -289 602 -282 630
rect -255 634 -250 643
rect -224 634 -219 643
rect -191 634 -186 643
rect -120 635 -115 644
rect -89 635 -84 644
rect -56 635 -51 644
rect -4 643 113 644
rect 10 642 113 643
rect -389 585 -385 590
rect -358 585 -354 590
rect -341 575 -336 598
rect -308 596 -282 602
rect -236 605 -231 629
rect -205 605 -200 629
rect -236 599 -186 605
rect -172 603 -167 629
rect -152 603 -148 627
rect -308 575 -303 596
rect -255 586 -249 591
rect -220 586 -218 591
rect -205 576 -200 599
rect -172 598 -148 603
rect -101 606 -96 630
rect -70 606 -65 630
rect -101 600 -51 606
rect -37 604 -32 630
rect -13 604 -8 632
rect 17 633 22 642
rect 48 633 53 642
rect 81 633 86 642
rect -172 597 -164 598
rect -172 576 -167 597
rect -118 587 -114 592
rect -85 587 -83 592
rect -70 577 -65 600
rect -37 598 -8 604
rect 36 604 41 628
rect 67 604 72 628
rect 36 598 86 604
rect 100 602 105 628
rect 116 602 123 712
rect 162 637 171 931
rect 513 1053 519 1235
rect 547 1226 551 1245
rect 576 1226 580 1245
rect 605 1226 609 1245
rect 634 1226 638 1245
rect 655 1231 696 1235
rect 655 1226 659 1231
rect 663 1226 667 1231
rect 692 1226 696 1231
rect 765 1226 769 1245
rect 794 1226 798 1245
rect 823 1226 827 1245
rect 852 1226 856 1245
rect 873 1231 914 1235
rect 873 1226 877 1231
rect 881 1226 885 1231
rect 910 1226 914 1231
rect 998 1228 1002 1246
rect 1027 1228 1031 1247
rect 1056 1228 1060 1247
rect 1085 1228 1089 1247
rect 1106 1233 1147 1237
rect 1106 1228 1110 1233
rect 1114 1228 1118 1233
rect 1143 1228 1147 1233
rect 1258 1229 1262 1248
rect 1287 1229 1291 1248
rect 1316 1229 1320 1248
rect 1345 1229 1349 1248
rect 1366 1234 1407 1238
rect 1366 1229 1370 1234
rect 1374 1229 1378 1234
rect 1403 1229 1407 1234
rect 548 1183 551 1188
rect 568 1154 572 1222
rect 575 1182 580 1187
rect 575 1166 578 1182
rect 597 1171 601 1222
rect 626 1215 630 1222
rect 655 1215 659 1222
rect 626 1212 659 1215
rect 684 1215 688 1222
rect 713 1215 717 1222
rect 684 1212 717 1215
rect 662 1193 670 1197
rect 667 1192 670 1193
rect 713 1189 717 1212
rect 713 1188 728 1189
rect 713 1179 719 1188
rect 768 1183 769 1188
rect 597 1166 699 1171
rect 597 1154 601 1166
rect 695 1165 699 1166
rect 713 1162 717 1179
rect 655 1154 659 1155
rect 713 1154 717 1157
rect 786 1154 790 1222
rect 793 1182 798 1187
rect 793 1167 796 1182
rect 815 1171 819 1222
rect 844 1215 848 1222
rect 873 1215 877 1222
rect 844 1212 877 1215
rect 902 1215 906 1222
rect 931 1215 935 1222
rect 902 1212 935 1215
rect 880 1193 888 1197
rect 885 1192 888 1193
rect 815 1166 917 1171
rect 815 1154 819 1166
rect 913 1165 917 1166
rect 931 1162 935 1212
rect 999 1185 1002 1190
rect 873 1154 877 1155
rect 931 1154 935 1157
rect 1019 1156 1023 1224
rect 1026 1189 1030 1190
rect 1026 1184 1031 1189
rect 1026 1175 1029 1184
rect 1048 1173 1052 1224
rect 1077 1217 1081 1224
rect 1106 1217 1110 1224
rect 1077 1214 1110 1217
rect 1135 1217 1139 1224
rect 1164 1217 1168 1224
rect 1135 1214 1168 1217
rect 1113 1195 1121 1199
rect 1118 1194 1121 1195
rect 1164 1191 1168 1214
rect 1164 1181 1200 1191
rect 1259 1186 1262 1191
rect 1048 1168 1150 1173
rect 1048 1156 1052 1168
rect 1146 1167 1150 1168
rect 1164 1164 1168 1181
rect 1106 1156 1110 1157
rect 1164 1156 1168 1159
rect 1279 1157 1283 1225
rect 1286 1185 1291 1190
rect 1286 1173 1289 1185
rect 1308 1174 1312 1225
rect 1337 1218 1341 1225
rect 1366 1218 1370 1225
rect 1337 1215 1370 1218
rect 1395 1218 1399 1225
rect 1424 1218 1428 1225
rect 1395 1215 1428 1218
rect 1373 1196 1381 1200
rect 1378 1195 1381 1196
rect 1424 1192 1428 1215
rect 1424 1191 1432 1192
rect 1424 1183 1473 1191
rect 1424 1182 1432 1183
rect 1308 1169 1410 1174
rect 1308 1157 1312 1169
rect 1406 1168 1410 1169
rect 1424 1165 1428 1182
rect 1366 1157 1370 1158
rect 1424 1157 1428 1160
rect 630 1150 634 1154
rect 688 1150 692 1154
rect 848 1150 852 1154
rect 906 1150 910 1154
rect 1081 1152 1085 1156
rect 1139 1152 1143 1156
rect 1341 1153 1345 1157
rect 1399 1153 1403 1157
rect 547 1146 551 1150
rect 576 1146 580 1150
rect 605 1146 609 1150
rect 663 1146 667 1150
rect 765 1146 769 1150
rect 794 1146 798 1150
rect 823 1146 827 1150
rect 881 1146 885 1150
rect 998 1148 1002 1152
rect 1027 1148 1031 1152
rect 1056 1148 1060 1152
rect 1114 1148 1118 1152
rect 995 1147 1183 1148
rect 944 1146 1253 1147
rect 1258 1146 1262 1153
rect 1287 1149 1291 1153
rect 1316 1149 1320 1153
rect 1374 1149 1378 1153
rect 1265 1148 1443 1149
rect 1265 1146 2990 1148
rect 544 1142 2990 1146
rect 544 1141 1274 1142
rect 1435 1141 2990 1142
rect 544 1140 999 1141
rect 544 1139 950 1140
rect 513 1047 783 1053
rect 1240 1050 1244 1051
rect 1139 1047 1409 1050
rect 513 1046 586 1047
rect 513 805 527 1046
rect 576 1028 580 1046
rect 605 1028 609 1047
rect 634 1028 638 1047
rect 663 1028 667 1047
rect 778 1044 783 1047
rect 1028 1044 1409 1047
rect 778 1043 1212 1044
rect 778 1038 1153 1043
rect 778 1037 1051 1038
rect 684 1033 725 1037
rect 684 1028 688 1033
rect 692 1028 696 1033
rect 721 1028 725 1033
rect 803 1028 808 1037
rect 834 1028 839 1037
rect 867 1028 872 1037
rect 597 1000 601 1024
rect 597 996 617 1000
rect 578 985 580 990
rect 597 956 601 996
rect 626 973 630 1024
rect 655 1017 659 1024
rect 684 1017 688 1024
rect 655 1014 688 1017
rect 713 1017 717 1024
rect 742 1017 746 1024
rect 713 1014 746 1017
rect 691 995 699 999
rect 696 994 699 995
rect 742 991 746 1014
rect 822 999 827 1023
rect 853 999 858 1023
rect 822 993 872 999
rect 742 988 750 991
rect 742 983 784 988
rect 742 981 750 983
rect 626 968 728 973
rect 626 956 630 968
rect 724 967 728 968
rect 742 964 746 981
rect 684 956 688 957
rect 742 956 746 959
rect 659 952 663 956
rect 717 952 721 956
rect 576 948 580 952
rect 605 948 609 952
rect 634 949 638 952
rect 632 948 638 949
rect 692 948 696 952
rect 548 941 754 948
rect 548 692 560 941
rect 777 846 784 983
rect 808 980 809 985
rect 839 980 840 985
rect 853 970 858 993
rect 886 970 891 1023
rect 1045 1014 1051 1037
rect 965 1009 1051 1014
rect 979 1003 983 1009
rect 1016 1003 1020 1009
rect 993 999 997 1003
rect 1007 979 1011 999
rect 1026 985 1030 999
rect 827 965 834 970
rect 960 972 982 976
rect 999 974 1000 978
rect 1007 975 1019 979
rect 1026 978 1029 985
rect 960 971 981 972
rect 803 961 808 965
rect 867 961 872 965
rect 797 960 898 961
rect 804 954 898 960
rect 812 898 941 905
rect 819 889 824 898
rect 850 889 855 898
rect 883 889 888 898
rect 838 860 843 884
rect 869 860 874 884
rect 838 854 888 860
rect 902 857 907 884
rect 960 857 967 971
rect 1007 970 1011 975
rect 989 967 1011 970
rect 989 962 993 967
rect 1007 962 1011 967
rect 1026 962 1030 978
rect 979 955 983 958
rect 997 955 1001 958
rect 1016 955 1020 958
rect 975 954 1039 955
rect 984 952 1039 954
rect 1044 905 1051 1009
rect 1007 898 1051 905
rect 777 841 825 846
rect 853 841 856 846
rect 588 792 768 798
rect 580 791 768 792
rect 586 772 590 791
rect 615 772 619 791
rect 644 772 648 791
rect 673 772 677 791
rect 694 777 735 781
rect 694 772 698 777
rect 702 772 706 777
rect 731 772 735 777
rect 587 729 590 734
rect 607 700 611 768
rect 636 717 640 768
rect 665 761 669 768
rect 694 761 698 768
rect 665 758 698 761
rect 723 761 727 768
rect 752 761 756 768
rect 723 758 756 761
rect 701 739 709 743
rect 706 738 709 739
rect 752 735 756 758
rect 752 725 760 735
rect 636 712 738 717
rect 636 700 640 712
rect 734 711 738 712
rect 752 708 756 725
rect 694 700 698 701
rect 752 700 756 703
rect 669 696 673 700
rect 727 696 731 700
rect 586 692 590 696
rect 615 692 619 696
rect 644 692 648 696
rect 702 692 706 696
rect 548 685 771 692
rect 548 637 560 685
rect 777 664 784 841
rect 869 831 874 854
rect 902 852 967 857
rect 902 831 907 852
rect 843 826 850 831
rect 819 822 824 826
rect 883 822 888 826
rect 621 657 784 664
rect 813 815 920 822
rect 162 630 560 637
rect 548 627 560 630
rect 813 627 827 815
rect 1139 802 1153 1038
rect 1202 1025 1206 1043
rect 1231 1025 1235 1044
rect 1260 1025 1264 1044
rect 1289 1025 1293 1044
rect 1404 1041 1409 1044
rect 1739 1044 2009 1050
rect 1739 1043 1812 1044
rect 1739 1042 1753 1043
rect 1672 1041 1753 1042
rect 1404 1034 1753 1041
rect 1310 1030 1351 1034
rect 1310 1025 1314 1030
rect 1318 1025 1322 1030
rect 1347 1025 1351 1030
rect 1429 1025 1434 1034
rect 1460 1025 1465 1034
rect 1493 1025 1498 1034
rect 1223 997 1227 1021
rect 1223 993 1243 997
rect 1204 982 1206 987
rect 1223 953 1227 993
rect 1252 970 1256 1021
rect 1281 1014 1285 1021
rect 1310 1014 1314 1021
rect 1281 1011 1314 1014
rect 1339 1014 1343 1021
rect 1368 1014 1372 1021
rect 1339 1011 1372 1014
rect 1317 992 1325 996
rect 1322 991 1325 992
rect 1368 988 1372 1011
rect 1448 996 1453 1020
rect 1479 996 1484 1020
rect 1448 990 1498 996
rect 1368 985 1376 988
rect 1368 980 1410 985
rect 1368 978 1376 980
rect 1252 965 1354 970
rect 1252 953 1256 965
rect 1350 964 1354 965
rect 1368 961 1372 978
rect 1310 953 1314 954
rect 1368 953 1372 956
rect 1285 949 1289 953
rect 1343 949 1347 953
rect 1202 945 1206 949
rect 1231 945 1235 949
rect 1260 945 1264 949
rect 1318 945 1322 949
rect 1174 938 1380 945
rect 548 624 827 627
rect 1174 689 1186 938
rect 1403 843 1410 980
rect 1434 977 1435 982
rect 1465 977 1466 982
rect 1479 967 1484 990
rect 1512 967 1517 1020
rect 1671 1011 1677 1034
rect 1591 1006 1677 1011
rect 1605 1000 1609 1006
rect 1642 1000 1646 1006
rect 1619 996 1623 1000
rect 1633 976 1637 996
rect 1652 979 1656 996
rect 1453 962 1460 967
rect 1586 969 1608 973
rect 1625 971 1626 975
rect 1633 972 1645 976
rect 1652 975 1659 979
rect 1586 968 1607 969
rect 1429 958 1434 962
rect 1493 958 1498 962
rect 1423 957 1524 958
rect 1430 951 1524 957
rect 1438 895 1567 902
rect 1445 886 1450 895
rect 1476 886 1481 895
rect 1509 886 1514 895
rect 1464 857 1469 881
rect 1495 857 1500 881
rect 1464 851 1514 857
rect 1528 854 1533 881
rect 1586 854 1593 968
rect 1633 967 1637 972
rect 1615 964 1637 967
rect 1615 959 1619 964
rect 1633 959 1637 964
rect 1652 959 1656 975
rect 1605 952 1609 955
rect 1623 952 1627 955
rect 1642 952 1646 955
rect 1601 951 1665 952
rect 1610 949 1665 951
rect 1670 902 1677 1006
rect 1633 895 1677 902
rect 1403 838 1451 843
rect 1479 838 1482 843
rect 1214 789 1394 795
rect 1206 788 1394 789
rect 1212 769 1216 788
rect 1241 769 1245 788
rect 1270 769 1274 788
rect 1299 769 1303 788
rect 1320 774 1361 778
rect 1320 769 1324 774
rect 1328 769 1332 774
rect 1357 769 1361 774
rect 1213 726 1216 731
rect 1233 697 1237 765
rect 1262 714 1266 765
rect 1291 758 1295 765
rect 1320 758 1324 765
rect 1291 755 1324 758
rect 1349 758 1353 765
rect 1378 758 1382 765
rect 1349 755 1382 758
rect 1327 736 1335 740
rect 1332 735 1335 736
rect 1378 732 1382 755
rect 1378 722 1386 732
rect 1262 709 1364 714
rect 1262 697 1266 709
rect 1360 708 1364 709
rect 1378 705 1382 722
rect 1320 697 1324 698
rect 1378 697 1382 700
rect 1295 693 1299 697
rect 1353 693 1357 697
rect 1212 689 1216 693
rect 1241 689 1245 693
rect 1270 689 1274 693
rect 1328 689 1332 693
rect 1174 682 1397 689
rect 1174 624 1186 682
rect 1403 661 1410 838
rect 1495 828 1500 851
rect 1528 849 1593 854
rect 1528 828 1533 849
rect 1469 823 1476 828
rect 1445 819 1450 823
rect 1509 819 1514 823
rect 1247 654 1410 661
rect 1439 812 1546 819
rect 1439 624 1453 812
rect 1739 802 1753 1034
rect 1802 1025 1806 1043
rect 1831 1025 1835 1044
rect 1839 1043 1843 1044
rect 1860 1025 1864 1044
rect 1889 1025 1893 1044
rect 2004 1041 2009 1044
rect 2342 1047 2612 1053
rect 2342 1046 2415 1047
rect 2004 1036 2277 1041
rect 2342 1036 2356 1046
rect 2004 1034 2356 1036
rect 1910 1030 1951 1034
rect 1910 1025 1914 1030
rect 1918 1025 1922 1030
rect 1947 1025 1951 1030
rect 2029 1025 2034 1034
rect 2060 1025 2065 1034
rect 2093 1025 2098 1034
rect 2271 1028 2356 1034
rect 1823 997 1827 1021
rect 1823 993 1843 997
rect 1804 982 1806 987
rect 1823 953 1827 993
rect 1852 970 1856 1021
rect 1881 1014 1885 1021
rect 1910 1014 1914 1021
rect 1881 1011 1914 1014
rect 1939 1014 1943 1021
rect 1968 1014 1972 1021
rect 1939 1011 1972 1014
rect 1917 992 1925 996
rect 1922 991 1925 992
rect 1968 988 1972 1011
rect 2048 996 2053 1020
rect 2079 996 2084 1020
rect 2048 990 2098 996
rect 1968 985 1976 988
rect 1968 980 2010 985
rect 1968 978 1976 980
rect 1852 965 1954 970
rect 1852 953 1856 965
rect 1950 964 1954 965
rect 1968 961 1972 978
rect 1910 953 1914 954
rect 1968 953 1972 956
rect 1885 949 1889 953
rect 1943 949 1947 953
rect 1802 945 1806 949
rect 1831 945 1835 949
rect 1860 945 1864 949
rect 1918 945 1922 949
rect 1774 938 1980 945
rect 548 620 1453 624
rect 1774 689 1786 938
rect 2003 843 2010 980
rect 2034 977 2035 982
rect 2065 977 2066 982
rect 2079 967 2084 990
rect 2112 967 2117 1020
rect 2271 1011 2277 1028
rect 2191 1006 2277 1011
rect 2205 1000 2209 1006
rect 2242 1000 2246 1006
rect 2219 996 2223 1000
rect 2233 976 2237 996
rect 2252 979 2256 996
rect 2053 962 2060 967
rect 2186 969 2208 973
rect 2225 971 2226 975
rect 2233 972 2245 976
rect 2252 975 2259 979
rect 2186 968 2207 969
rect 2029 958 2034 962
rect 2093 958 2098 962
rect 2023 957 2124 958
rect 2030 951 2124 957
rect 2038 895 2167 902
rect 2045 886 2050 895
rect 2076 886 2081 895
rect 2109 886 2114 895
rect 2064 857 2069 881
rect 2095 857 2100 881
rect 2064 851 2114 857
rect 2128 854 2133 881
rect 2186 854 2193 968
rect 2233 967 2237 972
rect 2215 964 2237 967
rect 2215 959 2219 964
rect 2233 959 2237 964
rect 2252 959 2256 975
rect 2205 952 2209 955
rect 2223 952 2227 955
rect 2242 952 2246 955
rect 2201 951 2265 952
rect 2210 949 2265 951
rect 2270 902 2277 1006
rect 2233 895 2277 902
rect 2003 838 2051 843
rect 2079 838 2082 843
rect 1814 789 1994 795
rect 1806 788 1994 789
rect 1812 769 1816 788
rect 1841 769 1845 788
rect 1870 769 1874 788
rect 1899 769 1903 788
rect 1920 774 1961 778
rect 1920 769 1924 774
rect 1928 769 1932 774
rect 1957 769 1961 774
rect 1814 726 1816 731
rect 1833 697 1837 765
rect 1862 714 1866 765
rect 1891 758 1895 765
rect 1920 758 1924 765
rect 1891 755 1924 758
rect 1949 758 1953 765
rect 1978 758 1982 765
rect 1949 755 1982 758
rect 1927 736 1935 740
rect 1932 735 1935 736
rect 1978 732 1982 755
rect 1978 722 1986 732
rect 1862 709 1964 714
rect 1862 697 1866 709
rect 1960 708 1964 709
rect 1978 705 1982 722
rect 1920 697 1924 698
rect 1978 697 1982 700
rect 1895 693 1899 697
rect 1953 693 1957 697
rect 1812 689 1816 693
rect 1841 689 1845 693
rect 1870 689 1874 693
rect 1928 689 1932 693
rect 1774 682 1997 689
rect 1774 624 1786 682
rect 2003 661 2010 838
rect 2095 828 2100 851
rect 2128 849 2193 854
rect 2128 828 2133 849
rect 2069 823 2076 828
rect 2045 819 2050 823
rect 2109 819 2114 823
rect 1847 654 2010 661
rect 2039 812 2146 819
rect 2039 624 2053 812
rect 2342 805 2356 1028
rect 2405 1028 2409 1046
rect 2434 1028 2438 1047
rect 2463 1028 2467 1047
rect 2492 1028 2496 1047
rect 2607 1044 2612 1047
rect 2607 1037 2880 1044
rect 2513 1033 2554 1037
rect 2513 1028 2517 1033
rect 2521 1028 2525 1033
rect 2550 1028 2554 1033
rect 2632 1028 2637 1037
rect 2663 1028 2668 1037
rect 2696 1028 2701 1037
rect 2426 1000 2430 1024
rect 2426 996 2446 1000
rect 2407 985 2409 990
rect 2426 956 2430 996
rect 2455 973 2459 1024
rect 2484 1017 2488 1024
rect 2513 1017 2517 1024
rect 2484 1014 2517 1017
rect 2542 1017 2546 1024
rect 2571 1017 2575 1024
rect 2542 1014 2575 1017
rect 2520 995 2528 999
rect 2525 994 2528 995
rect 2571 991 2575 1014
rect 2651 999 2656 1023
rect 2682 999 2687 1023
rect 2651 993 2701 999
rect 2571 988 2579 991
rect 2571 983 2613 988
rect 2571 981 2579 983
rect 2455 968 2557 973
rect 2455 956 2459 968
rect 2553 967 2557 968
rect 2571 964 2575 981
rect 2513 956 2517 957
rect 2571 956 2575 959
rect 2488 952 2492 956
rect 2546 952 2550 956
rect 2405 948 2409 952
rect 2434 948 2438 952
rect 2463 950 2467 952
rect 2462 948 2467 950
rect 2521 948 2525 952
rect 2377 941 2583 948
rect 1774 623 2053 624
rect 2377 692 2389 941
rect 2606 846 2613 983
rect 2637 980 2638 985
rect 2668 980 2669 985
rect 2682 970 2687 993
rect 2715 970 2720 1023
rect 2874 1014 2880 1037
rect 2794 1009 2880 1014
rect 2808 1003 2812 1009
rect 2845 1003 2849 1009
rect 2822 999 2826 1003
rect 2836 979 2840 999
rect 2855 982 2859 999
rect 2656 965 2663 970
rect 2789 972 2811 976
rect 2828 974 2829 978
rect 2836 975 2848 979
rect 2855 978 2864 982
rect 2789 971 2810 972
rect 2632 961 2637 965
rect 2696 961 2701 965
rect 2626 960 2727 961
rect 2633 954 2727 960
rect 2641 898 2770 905
rect 2648 889 2653 898
rect 2679 889 2684 898
rect 2712 889 2717 898
rect 2667 860 2672 884
rect 2698 860 2703 884
rect 2667 854 2717 860
rect 2731 857 2736 884
rect 2789 857 2796 971
rect 2836 970 2840 975
rect 2818 967 2840 970
rect 2818 962 2822 967
rect 2836 962 2840 967
rect 2855 962 2859 978
rect 2808 955 2812 958
rect 2826 955 2830 958
rect 2845 955 2849 958
rect 2804 954 2868 955
rect 2813 952 2868 954
rect 2873 905 2880 1009
rect 2836 898 2880 905
rect 2606 841 2654 846
rect 2682 841 2685 846
rect 2417 792 2597 798
rect 2409 791 2597 792
rect 2415 772 2419 791
rect 2444 772 2448 791
rect 2473 772 2477 791
rect 2502 772 2506 791
rect 2523 777 2564 781
rect 2523 772 2527 777
rect 2531 772 2535 777
rect 2560 772 2564 777
rect 2416 729 2419 734
rect 2436 700 2440 768
rect 2465 717 2469 768
rect 2494 761 2498 768
rect 2523 761 2527 768
rect 2494 758 2527 761
rect 2552 761 2556 768
rect 2581 761 2585 768
rect 2552 758 2585 761
rect 2530 739 2538 743
rect 2535 738 2538 739
rect 2581 735 2585 758
rect 2581 725 2589 735
rect 2465 712 2567 717
rect 2465 700 2469 712
rect 2563 711 2567 712
rect 2581 708 2585 725
rect 2523 700 2527 701
rect 2581 700 2585 703
rect 2498 696 2502 700
rect 2556 696 2560 700
rect 2415 692 2419 696
rect 2444 692 2448 696
rect 2473 692 2477 696
rect 2531 692 2535 696
rect 2377 685 2600 692
rect 2377 627 2389 685
rect 2606 664 2613 841
rect 2698 831 2703 854
rect 2731 852 2796 857
rect 2731 831 2736 852
rect 2672 826 2679 831
rect 2648 822 2653 826
rect 2712 822 2717 826
rect 2450 657 2613 664
rect 2642 815 2749 822
rect 2642 627 2656 815
rect 2377 625 2656 627
rect 2971 625 2989 1141
rect 2377 623 2989 625
rect 1774 620 2989 623
rect 548 619 2989 620
rect 548 618 827 619
rect 1174 618 2989 619
rect 1174 615 2053 618
rect 2630 617 2989 618
rect -37 577 -32 598
rect 18 585 23 590
rect 52 585 54 590
rect -367 570 -360 575
rect -231 571 -224 576
rect -96 572 -89 577
rect 67 575 72 598
rect 100 596 123 602
rect 100 575 105 596
rect -391 566 -386 570
rect -327 566 -322 570
rect -255 567 -250 571
rect -191 567 -186 571
rect -120 568 -115 572
rect -56 568 -51 572
rect 41 570 48 575
rect -261 566 -148 567
rect -126 566 -13 568
rect 17 566 22 570
rect 81 566 86 570
rect -397 565 -284 566
rect -261 565 149 566
rect -397 564 149 565
rect -398 561 149 564
rect -397 560 -141 561
rect -397 559 -284 560
rect 11 559 149 561
rect -123 532 -20 533
rect -154 530 121 532
rect -423 527 -296 529
rect -253 527 121 530
rect -423 526 121 527
rect -423 524 -150 526
rect -423 522 -296 524
rect -253 523 -150 524
rect -392 513 -387 522
rect -361 513 -356 522
rect -328 513 -323 522
rect -246 514 -241 523
rect -215 514 -210 523
rect -182 514 -177 523
rect -116 517 -111 526
rect -85 517 -80 526
rect -52 517 -47 526
rect 18 525 121 526
rect -373 484 -368 508
rect -342 484 -337 508
rect -373 478 -323 484
rect -309 482 -304 508
rect -227 485 -222 509
rect -196 485 -191 509
rect -392 465 -386 470
rect -357 465 -355 470
rect -342 455 -337 478
rect -309 476 -303 482
rect -227 479 -177 485
rect -163 482 -158 509
rect -97 488 -92 512
rect -66 488 -61 512
rect -97 482 -47 488
rect -33 486 -28 512
rect 25 516 30 525
rect 56 516 61 525
rect 89 516 94 525
rect 44 487 49 511
rect 75 487 80 511
rect -309 455 -304 476
rect -245 466 -240 471
rect -212 466 -209 471
rect -196 456 -191 479
rect -163 476 -155 482
rect -163 456 -158 476
rect -116 469 -110 474
rect -83 469 -79 474
rect -66 459 -61 482
rect -33 480 -25 486
rect 44 481 94 487
rect 108 485 113 511
rect -33 459 -28 480
rect 25 468 31 473
rect 58 468 62 473
rect -368 450 -361 455
rect -222 451 -215 456
rect -92 454 -85 459
rect 75 458 80 481
rect 108 479 115 485
rect 108 458 113 479
rect -392 446 -387 450
rect -328 446 -323 450
rect -246 447 -241 451
rect -182 447 -177 451
rect -116 450 -111 454
rect -52 450 -47 454
rect 49 453 56 458
rect -122 448 -9 450
rect 25 449 30 453
rect 89 449 94 453
rect 141 449 149 559
rect -152 447 -9 448
rect 19 447 149 449
rect -291 446 149 447
rect -413 445 149 446
rect -503 444 149 445
rect -503 443 -9 444
rect -503 441 -118 443
rect 19 442 149 444
rect -413 440 -118 441
rect -413 439 -251 440
rect -890 321 -540 326
rect -1054 268 -921 274
rect -1047 259 -1042 268
rect -1016 259 -1011 268
rect -983 259 -978 268
rect -1028 230 -1023 254
rect -997 230 -992 254
rect -1096 223 -1054 226
rect -1028 224 -978 230
rect -964 225 -959 254
rect -1057 216 -1054 223
rect -1057 211 -1041 216
rect -997 201 -992 224
rect -964 201 -959 218
rect -1023 196 -1016 201
rect -1047 192 -1042 196
rect -983 192 -978 196
rect -1278 117 -1274 186
rect -1193 183 -1111 189
rect -1053 185 -955 192
rect -1193 173 -1189 183
rect -1116 173 -1013 176
rect -1241 144 -1237 169
rect -1260 143 -1162 144
rect -1260 134 -1174 143
rect -1163 134 -1162 143
rect -1116 117 -1111 173
rect -929 166 -921 268
rect -881 218 -798 225
rect -1052 160 -921 166
rect -1045 151 -1040 160
rect -1014 151 -1009 160
rect -981 151 -976 160
rect -1278 112 -1111 117
rect -1026 122 -1021 146
rect -995 122 -990 146
rect -1026 116 -976 122
rect -1043 103 -1039 108
rect -1008 108 -1004 109
rect -1008 102 -1004 103
rect -995 93 -990 116
rect -962 115 -957 146
rect -804 148 -798 218
rect -645 177 -639 262
rect -114 225 -11 226
rect 1907 225 2423 226
rect -411 224 -276 225
rect -266 224 -124 225
rect -114 224 14 225
rect 1169 224 2423 225
rect -411 223 2423 224
rect -557 220 2423 223
rect -548 219 2423 220
rect -548 218 -146 219
rect -548 213 -404 218
rect -385 217 -282 218
rect -804 140 -498 148
rect -962 111 -893 115
rect -962 93 -957 111
rect -1021 88 -1014 93
rect -1045 84 -1040 88
rect -981 84 -976 88
rect -1051 77 -953 84
rect -896 -300 -893 111
rect -410 104 -405 213
rect -378 208 -373 217
rect -347 208 -342 217
rect -314 208 -309 217
rect -242 209 -237 218
rect -211 209 -206 218
rect -178 209 -173 218
rect -107 210 -102 219
rect -76 210 -71 219
rect -43 210 -38 219
rect 9 218 2423 219
rect 23 217 126 218
rect -359 179 -354 203
rect -328 179 -323 203
rect -359 173 -309 179
rect -295 177 -290 203
rect -223 180 -218 204
rect -192 180 -187 204
rect -376 160 -372 165
rect -345 160 -341 165
rect -328 150 -323 173
rect -295 171 -285 177
rect -295 150 -290 171
rect -223 174 -173 180
rect -159 178 -154 204
rect -88 181 -83 205
rect -57 181 -52 205
rect -241 161 -236 166
rect -207 161 -205 166
rect -192 151 -187 174
rect -159 172 -146 178
rect -159 151 -154 172
rect -88 175 -38 181
rect -24 179 -19 205
rect 30 208 35 217
rect 61 208 66 217
rect 94 208 99 217
rect -106 162 -101 167
rect -72 162 -70 167
rect -57 152 -52 175
rect -24 173 -9 179
rect -24 152 -19 173
rect 49 179 54 203
rect 80 179 85 203
rect 49 173 99 179
rect 113 177 118 203
rect 32 160 36 165
rect 65 160 67 165
rect -354 145 -347 150
rect -218 146 -211 151
rect -83 147 -76 152
rect 80 150 85 173
rect 113 171 1785 177
rect 113 150 118 171
rect -378 141 -373 145
rect -314 141 -309 145
rect -242 142 -237 146
rect -178 142 -173 146
rect -107 143 -102 147
rect -43 143 -38 147
rect 54 145 61 150
rect -248 141 -135 142
rect -113 141 0 143
rect 30 141 35 145
rect 94 141 99 145
rect -384 140 -271 141
rect -248 140 162 141
rect -384 139 162 140
rect -385 136 162 139
rect -384 135 -128 136
rect -384 134 -271 135
rect 24 134 162 136
rect -110 107 -7 108
rect -141 105 134 107
rect -410 102 -283 104
rect -240 102 134 105
rect -410 101 134 102
rect -410 99 -137 101
rect -410 97 -283 99
rect -240 98 -137 99
rect -379 88 -374 97
rect -348 88 -343 97
rect -315 88 -310 97
rect -233 89 -228 98
rect -202 89 -197 98
rect -169 89 -164 98
rect -103 92 -98 101
rect -72 92 -67 101
rect -39 92 -34 101
rect 31 100 134 101
rect -360 59 -355 83
rect -329 59 -324 83
rect -360 53 -310 59
rect -296 58 -291 83
rect -214 60 -209 84
rect -183 60 -178 84
rect -296 57 -281 58
rect -378 40 -373 45
rect -344 40 -342 45
rect -329 30 -324 53
rect -296 50 -283 57
rect -214 54 -164 60
rect -150 57 -145 84
rect -84 63 -79 87
rect -53 63 -48 87
rect -84 57 -34 63
rect -20 61 -15 87
rect 38 91 43 100
rect 69 91 74 100
rect 102 91 107 100
rect 57 62 62 86
rect 88 62 93 86
rect -296 30 -291 50
rect -231 41 -227 46
rect -199 41 -196 46
rect -183 31 -178 54
rect -150 51 -140 57
rect -150 31 -145 51
rect -102 44 -97 49
rect -70 44 -66 49
rect -53 34 -48 57
rect -20 55 -8 61
rect 57 56 107 62
rect 121 60 126 86
rect -20 34 -15 55
rect 40 43 44 48
rect 71 43 75 48
rect -355 25 -348 30
rect -209 26 -202 31
rect -79 29 -72 34
rect 88 33 93 56
rect 121 54 132 60
rect 121 33 126 54
rect -645 21 -396 22
rect -379 21 -374 25
rect -315 21 -310 25
rect -233 22 -228 26
rect -169 22 -164 26
rect -103 25 -98 29
rect -39 25 -34 29
rect 62 28 69 33
rect -109 23 -4 25
rect 38 24 43 28
rect 102 24 107 28
rect 154 24 162 134
rect 32 23 135 24
rect -125 22 135 23
rect -263 21 135 22
rect 146 21 162 24
rect -645 20 -281 21
rect -263 20 162 21
rect -645 18 162 20
rect -645 17 -85 18
rect 32 17 162 18
rect -645 16 -139 17
rect -636 15 -139 16
rect -125 15 -105 17
rect -636 14 -281 15
rect -263 14 -238 15
rect -636 9 -396 14
rect -666 -225 -353 -224
rect -666 -226 -94 -225
rect -62 -226 41 -224
rect -666 -231 178 -226
rect -666 -232 -94 -231
rect -666 -234 -353 -232
rect -333 -233 -230 -232
rect -896 -310 -446 -300
rect -358 -346 -353 -234
rect -326 -242 -321 -233
rect -295 -242 -290 -233
rect -262 -242 -257 -233
rect -190 -241 -185 -232
rect -159 -241 -154 -232
rect -126 -241 -121 -232
rect -55 -240 -50 -231
rect -24 -240 -19 -231
rect 9 -240 14 -231
rect 61 -232 178 -231
rect 75 -233 178 -232
rect -307 -271 -302 -247
rect -276 -271 -271 -247
rect -307 -277 -257 -271
rect -243 -273 -238 -247
rect -171 -270 -166 -246
rect -140 -270 -135 -246
rect -323 -290 -320 -285
rect -293 -290 -289 -285
rect -276 -300 -271 -277
rect -243 -280 -229 -273
rect -171 -276 -121 -270
rect -107 -272 -102 -246
rect -36 -269 -31 -245
rect -5 -269 0 -245
rect -243 -300 -238 -280
rect -187 -288 -184 -284
rect -193 -289 -184 -288
rect -155 -289 -153 -284
rect -140 -299 -135 -276
rect -107 -278 -74 -272
rect -36 -275 14 -269
rect 28 -271 33 -245
rect 82 -242 87 -233
rect 113 -242 118 -233
rect 146 -242 151 -233
rect 101 -271 106 -247
rect 132 -271 137 -247
rect -107 -299 -102 -278
rect -55 -288 -49 -283
rect -20 -288 -18 -283
rect -5 -298 0 -275
rect 28 -277 62 -271
rect 101 -277 151 -271
rect 165 -272 170 -247
rect 28 -298 33 -277
rect 79 -290 82 -285
rect 87 -290 88 -285
rect 117 -290 119 -285
rect -302 -305 -295 -300
rect -166 -304 -159 -299
rect -31 -303 -24 -298
rect 132 -300 137 -277
rect 165 -280 345 -272
rect 165 -300 170 -280
rect -326 -309 -321 -305
rect -262 -309 -257 -305
rect -190 -308 -185 -304
rect -126 -308 -121 -304
rect -55 -307 -50 -303
rect 9 -307 14 -303
rect 106 -305 113 -300
rect -196 -309 -83 -308
rect -61 -309 52 -307
rect 82 -309 87 -305
rect 146 -309 151 -305
rect -332 -310 -219 -309
rect -196 -310 214 -309
rect -332 -311 214 -310
rect -333 -314 214 -311
rect -332 -315 -76 -314
rect -332 -316 -219 -315
rect 76 -316 214 -314
rect -58 -343 45 -342
rect -89 -345 175 -343
rect -358 -348 -231 -346
rect -188 -348 175 -345
rect -358 -349 175 -348
rect -358 -351 -85 -349
rect -358 -353 -231 -351
rect -188 -352 -85 -351
rect -327 -362 -322 -353
rect -296 -362 -291 -353
rect -263 -362 -258 -353
rect -181 -361 -176 -352
rect -150 -361 -145 -352
rect -117 -361 -112 -352
rect -51 -358 -46 -349
rect -20 -358 -15 -349
rect 13 -358 18 -349
rect 83 -350 186 -349
rect -308 -391 -303 -367
rect -277 -391 -272 -367
rect -308 -397 -258 -391
rect -244 -393 -239 -367
rect -162 -390 -157 -366
rect -131 -390 -126 -366
rect -823 -406 -746 -404
rect -721 -406 -321 -405
rect -823 -410 -321 -406
rect -292 -410 -290 -405
rect -823 -411 -700 -410
rect -823 -413 -746 -411
rect -277 -420 -272 -397
rect -244 -399 -200 -393
rect -162 -396 -112 -390
rect -98 -393 -93 -366
rect -32 -387 -27 -363
rect -1 -387 4 -363
rect -32 -393 18 -387
rect 32 -389 37 -363
rect 90 -359 95 -350
rect 121 -359 126 -350
rect 154 -359 159 -350
rect 109 -388 114 -364
rect 140 -388 145 -364
rect -244 -420 -239 -399
rect -303 -425 -296 -420
rect -203 -417 -200 -399
rect -181 -409 -175 -404
rect -147 -409 -144 -404
rect -131 -419 -126 -396
rect -98 -399 -92 -393
rect -98 -419 -93 -399
rect -49 -406 -45 -401
rect -18 -406 -14 -401
rect -1 -416 4 -393
rect 32 -395 47 -389
rect 109 -394 159 -388
rect 173 -390 178 -364
rect 173 -391 180 -390
rect 32 -416 37 -395
rect 93 -407 96 -402
rect 123 -407 127 -402
rect -157 -424 -150 -419
rect -27 -421 -20 -416
rect 140 -417 145 -394
rect 173 -396 179 -391
rect 173 -417 178 -396
rect -327 -429 -322 -425
rect -263 -429 -258 -425
rect -181 -428 -176 -424
rect -117 -428 -112 -424
rect -51 -425 -46 -421
rect 13 -425 18 -421
rect 114 -422 121 -417
rect -57 -427 56 -425
rect 90 -426 95 -422
rect 154 -426 159 -422
rect 206 -426 214 -316
rect -87 -428 56 -427
rect 84 -428 214 -426
rect -226 -429 214 -428
rect -348 -430 214 -429
rect -634 -431 214 -430
rect -634 -432 56 -431
rect -634 -435 -53 -432
rect 84 -433 214 -431
rect -634 -436 -186 -435
rect -634 -438 -346 -436
rect -571 -1574 -554 -438
rect -383 -595 -377 -438
rect -226 -499 -221 -444
rect -292 -503 -221 -499
rect -201 -499 -197 -444
rect -292 -571 -289 -503
rect -201 -504 -163 -499
rect -277 -518 -179 -512
rect -277 -519 -174 -518
rect -270 -528 -265 -519
rect -239 -528 -234 -519
rect -206 -528 -201 -519
rect -251 -557 -246 -533
rect -220 -557 -215 -533
rect -251 -563 -201 -557
rect -187 -560 -182 -533
rect -292 -576 -264 -571
rect -235 -575 -233 -571
rect -220 -586 -215 -563
rect -187 -565 -179 -560
rect -187 -586 -182 -565
rect -167 -576 -163 -504
rect -72 -543 -69 -444
rect 340 -465 345 -280
rect 1775 -305 1781 171
rect 2016 52 2174 58
rect 1799 2 2000 5
rect 2016 -296 2023 52
rect 2059 35 2155 36
rect 2059 34 2145 35
rect 2033 27 2145 34
rect 2033 -159 2042 27
rect 2059 26 2155 27
rect 2077 14 2081 26
rect 2089 -11 2095 -7
rect 2125 -8 2129 10
rect 2170 -8 2174 52
rect 2089 -12 2094 -11
rect 2059 -16 2094 -12
rect 2125 -14 2174 -8
rect 2289 -13 2294 168
rect 2415 32 2422 218
rect 2584 34 2680 37
rect 2852 34 2948 37
rect 2584 32 2948 34
rect 2415 31 2948 32
rect 2337 29 2948 31
rect 2337 28 2680 29
rect 2337 23 2425 28
rect 2584 27 2680 28
rect 2852 27 2948 29
rect 2329 21 2425 23
rect 2347 9 2351 21
rect 2602 15 2606 27
rect 2870 15 2874 27
rect 2359 -13 2365 -12
rect 2125 -24 2129 -14
rect 2289 -16 2365 -13
rect 2395 -13 2399 5
rect 2602 -10 2620 -6
rect 2650 -7 2654 11
rect 2650 -13 2698 -7
rect 2886 -10 2888 -6
rect 2918 -7 2922 11
rect 2395 -19 2398 -13
rect 2077 -53 2081 -28
rect 2395 -29 2399 -19
rect 2650 -23 2654 -13
rect 2918 -14 2921 -7
rect 2918 -23 2922 -14
rect 2058 -58 2136 -53
rect 2148 -58 2155 -53
rect 2347 -58 2351 -33
rect 2602 -52 2606 -27
rect 2870 -52 2874 -27
rect 2583 -56 2948 -52
rect 2583 -57 2680 -56
rect 2422 -58 2680 -57
rect 2851 -58 2948 -56
rect 2058 -59 2155 -58
rect 2328 -59 2605 -58
rect 2151 -61 2605 -59
rect 2151 -63 2425 -61
rect 2328 -64 2425 -63
rect 3229 -62 3235 -55
rect 3229 -67 3427 -62
rect 3229 -156 3235 -67
rect 3423 -110 3428 -67
rect 3414 -118 3600 -110
rect 3426 -133 3430 -118
rect 3559 -133 3563 -118
rect 3455 -137 3460 -133
rect 3489 -137 3493 -133
rect 3522 -137 3526 -133
rect 2212 -157 2502 -156
rect 2212 -158 2504 -157
rect 2594 -158 3252 -156
rect 2212 -159 3252 -158
rect 2033 -161 3252 -159
rect 2033 -163 2883 -161
rect 2033 -164 2504 -163
rect 2033 -238 2042 -164
rect 2212 -170 2504 -164
rect 2212 -171 2488 -170
rect 2219 -183 2223 -171
rect 2263 -183 2267 -171
rect 2307 -183 2311 -171
rect 2351 -183 2355 -171
rect 2395 -183 2399 -171
rect 2439 -183 2443 -171
rect 2255 -198 2259 -187
rect 2299 -198 2303 -187
rect 2343 -198 2347 -187
rect 2387 -198 2391 -187
rect 2431 -198 2435 -187
rect 2255 -202 2435 -198
rect 2431 -236 2440 -202
rect 2475 -233 2479 -187
rect 2494 -215 2504 -170
rect 2594 -170 2883 -163
rect 2890 -164 3252 -161
rect 2890 -170 2891 -164
rect 2594 -171 2870 -170
rect 2976 -171 3252 -164
rect 2601 -183 2605 -171
rect 2645 -183 2649 -171
rect 2689 -183 2693 -171
rect 2733 -183 2737 -171
rect 2777 -183 2781 -171
rect 2821 -183 2825 -171
rect 2983 -183 2987 -171
rect 3027 -183 3031 -171
rect 3071 -183 3075 -171
rect 3115 -183 3119 -171
rect 3159 -183 3163 -171
rect 3203 -183 3207 -171
rect 3405 -178 3411 -177
rect 3430 -178 3434 -177
rect 3405 -183 3434 -178
rect 3467 -182 3469 -178
rect 2637 -198 2641 -187
rect 2681 -198 2685 -187
rect 2725 -198 2729 -187
rect 2769 -198 2773 -187
rect 2813 -198 2817 -187
rect 2637 -202 2817 -198
rect 2475 -234 2487 -233
rect 2033 -245 2137 -238
rect 2041 -254 2046 -245
rect 2072 -254 2077 -245
rect 2105 -254 2110 -245
rect 2214 -249 2226 -240
rect 2262 -250 2271 -241
rect 2310 -251 2319 -242
rect 2356 -251 2362 -242
rect 2060 -283 2065 -259
rect 2091 -283 2096 -259
rect 2060 -289 2110 -283
rect 2124 -286 2129 -259
rect 2310 -278 2313 -251
rect 2403 -253 2406 -244
rect 2431 -245 2447 -236
rect 2431 -286 2435 -245
rect 2475 -286 2479 -234
rect 2486 -245 2487 -234
rect 2813 -236 2822 -202
rect 2857 -233 2861 -187
rect 3019 -198 3023 -187
rect 3063 -198 3067 -187
rect 3107 -198 3111 -187
rect 3151 -198 3155 -187
rect 3195 -198 3199 -187
rect 3019 -202 3199 -198
rect 2857 -234 2869 -233
rect 2599 -242 2608 -240
rect 2604 -248 2608 -242
rect 2599 -249 2608 -248
rect 2644 -243 2653 -241
rect 2649 -249 2653 -243
rect 2644 -250 2653 -249
rect 2695 -251 2701 -242
rect 2735 -251 2744 -242
rect 2779 -245 2788 -244
rect 2735 -271 2740 -251
rect 2783 -252 2788 -245
rect 2779 -253 2788 -252
rect 2813 -245 2829 -236
rect 2857 -245 2864 -234
rect 3195 -236 3204 -202
rect 3239 -233 3243 -187
rect 3239 -234 3251 -233
rect 2813 -286 2817 -245
rect 2857 -286 2861 -245
rect 2987 -249 2990 -240
rect 3031 -250 3035 -241
rect 3080 -251 3083 -242
rect 3123 -251 3126 -242
rect 3157 -244 3166 -243
rect 3157 -253 3170 -244
rect 3195 -245 3211 -236
rect 3239 -244 3245 -234
rect 3239 -245 3251 -244
rect 3157 -271 3162 -253
rect 3195 -286 3199 -245
rect 3239 -286 3243 -245
rect 2016 -297 2042 -296
rect 2070 -297 2074 -296
rect 2016 -302 2047 -297
rect 2070 -302 2078 -297
rect 2070 -305 2074 -302
rect 1775 -309 2074 -305
rect 1775 -310 1781 -309
rect 2091 -312 2096 -289
rect 2124 -292 2166 -286
rect 2259 -290 2263 -286
rect 2303 -290 2307 -286
rect 2347 -290 2351 -286
rect 2391 -290 2395 -286
rect 2641 -290 2645 -286
rect 2685 -290 2689 -286
rect 2729 -290 2733 -286
rect 2773 -290 2777 -286
rect 3023 -290 3027 -286
rect 3067 -290 3071 -286
rect 3111 -290 3115 -286
rect 3155 -290 3159 -286
rect 2124 -312 2129 -292
rect 2065 -317 2072 -312
rect 2041 -321 2046 -317
rect 2105 -321 2110 -317
rect 2035 -322 2137 -321
rect 2043 -328 2137 -322
rect 2162 -386 2165 -292
rect 2176 -309 2177 -306
rect 2219 -304 2223 -290
rect 2439 -304 2443 -290
rect 2601 -304 2605 -290
rect 2821 -304 2825 -290
rect 2983 -304 2987 -290
rect 3203 -304 3207 -290
rect 2216 -306 2492 -304
rect 2182 -309 2492 -306
rect 2216 -315 2492 -309
rect 2598 -313 2874 -304
rect 2980 -313 3256 -304
rect 2598 -315 3256 -313
rect 2216 -317 3256 -315
rect 2216 -319 2874 -317
rect 2980 -319 3256 -317
rect 3405 -386 3411 -183
rect 3551 -178 3555 -137
rect 3584 -178 3588 -137
rect 3498 -179 3501 -178
rect 3498 -183 3502 -179
rect 3498 -184 3501 -183
rect 3533 -184 3535 -180
rect 3551 -182 3567 -178
rect 3584 -182 3597 -178
rect 3551 -194 3555 -182
rect 3451 -198 3555 -194
rect 3451 -215 3455 -198
rect 3485 -215 3489 -198
rect 3518 -215 3522 -198
rect 3551 -215 3555 -198
rect 3584 -215 3588 -182
rect 3426 -227 3430 -219
rect 3460 -227 3464 -219
rect 3493 -227 3497 -219
rect 3526 -227 3530 -219
rect 3559 -227 3563 -219
rect 3423 -235 3607 -227
rect 2162 -387 2192 -386
rect 2205 -387 3411 -386
rect 2162 -391 3411 -387
rect 2162 -392 2192 -391
rect 2205 -392 3411 -391
rect 398 -413 497 -406
rect 401 -422 406 -413
rect 432 -422 437 -413
rect 465 -422 470 -413
rect 420 -451 425 -427
rect 451 -451 456 -427
rect 420 -457 470 -451
rect 484 -454 489 -427
rect 2287 -435 2819 -434
rect 2210 -440 2819 -435
rect 340 -469 407 -465
rect 401 -470 407 -469
rect 437 -470 438 -465
rect 451 -480 456 -457
rect 484 -459 492 -454
rect 484 -480 489 -459
rect 2039 -466 2203 -465
rect 425 -485 432 -480
rect 401 -489 406 -485
rect 465 -489 470 -485
rect 395 -496 502 -489
rect -73 -556 -69 -543
rect -101 -557 -69 -556
rect -111 -560 -69 -557
rect -246 -591 -239 -586
rect -270 -595 -265 -591
rect -206 -595 -201 -591
rect -383 -602 -169 -595
rect -189 -652 -182 -602
rect -111 -628 -106 -560
rect -101 -574 -11 -568
rect -5 -574 2 -568
rect -101 -575 2 -574
rect -94 -584 -89 -575
rect -63 -584 -58 -575
rect -30 -584 -25 -575
rect 153 -584 212 -578
rect 220 -584 256 -578
rect 153 -585 256 -584
rect -75 -613 -70 -589
rect -44 -613 -39 -589
rect -75 -619 -25 -613
rect -11 -616 -6 -589
rect 160 -594 165 -585
rect 191 -594 196 -585
rect 224 -594 229 -585
rect -94 -628 -88 -627
rect -111 -632 -88 -628
rect -59 -632 -57 -627
rect -44 -642 -39 -619
rect -11 -621 -3 -616
rect -11 -642 -6 -621
rect 179 -623 184 -599
rect 210 -623 215 -599
rect 179 -629 229 -623
rect 243 -626 248 -599
rect 163 -642 166 -637
rect 195 -642 197 -637
rect -70 -647 -63 -642
rect -94 -651 -89 -647
rect -30 -651 -25 -647
rect -100 -652 7 -651
rect 210 -652 215 -629
rect 243 -631 251 -626
rect 243 -652 248 -631
rect -189 -658 7 -652
rect 184 -657 191 -652
rect -2 -664 6 -658
rect 160 -661 165 -657
rect 224 -661 229 -657
rect 154 -663 261 -661
rect 462 -663 469 -496
rect 154 -664 469 -663
rect -1 -668 469 -664
rect -1 -669 160 -668
rect 462 -669 469 -668
rect 1976 -712 1983 -466
rect 1992 -477 2462 -466
rect 2057 -510 2061 -477
rect 2091 -510 2095 -477
rect 2124 -510 2128 -477
rect 2156 -510 2160 -477
rect 2179 -478 2462 -477
rect 2211 -491 2275 -485
rect 2211 -510 2215 -491
rect 2243 -510 2247 -491
rect 2058 -554 2060 -548
rect 2003 -570 2032 -567
rect 2080 -599 2084 -514
rect 2114 -549 2118 -514
rect 2147 -538 2151 -514
rect 2179 -538 2183 -514
rect 2188 -538 2192 -514
rect 2220 -538 2224 -514
rect 2271 -535 2275 -491
rect 2147 -542 2224 -538
rect 2270 -540 2387 -535
rect 2089 -555 2096 -549
rect 2114 -555 2163 -549
rect 2089 -565 2092 -555
rect 2114 -599 2118 -555
rect 2223 -579 2227 -574
rect 2271 -584 2275 -540
rect 2179 -588 2275 -584
rect 2179 -599 2183 -588
rect 2243 -599 2247 -588
rect 2151 -603 2156 -599
rect 2215 -603 2220 -599
rect 2057 -620 2061 -603
rect 2091 -620 2095 -603
rect 2124 -620 2128 -603
rect 2188 -620 2192 -603
rect 2050 -635 2207 -620
rect 1976 -723 2202 -712
rect 1976 -938 1983 -723
rect 2038 -724 2202 -723
rect 2056 -757 2060 -724
rect 2090 -757 2094 -724
rect 2123 -757 2127 -724
rect 2155 -757 2159 -724
rect 2210 -738 2275 -732
rect 2210 -757 2214 -738
rect 2242 -757 2246 -738
rect 2055 -801 2059 -795
rect 2005 -816 2039 -810
rect 2079 -846 2083 -761
rect 2113 -796 2117 -761
rect 2146 -785 2150 -761
rect 2178 -785 2182 -761
rect 2187 -785 2191 -761
rect 2219 -785 2223 -761
rect 2146 -789 2223 -785
rect 2088 -802 2095 -796
rect 2113 -802 2162 -796
rect 2089 -811 2092 -802
rect 2113 -846 2117 -802
rect 2270 -809 2275 -738
rect 2314 -809 2325 -664
rect 2362 -809 2369 -808
rect 2269 -814 2369 -809
rect 2222 -826 2226 -821
rect 2270 -831 2275 -814
rect 2314 -815 2325 -814
rect 2178 -835 2275 -831
rect 2362 -834 2369 -814
rect 2178 -846 2182 -835
rect 2242 -846 2246 -835
rect 2150 -850 2155 -846
rect 2214 -850 2219 -846
rect 2056 -867 2060 -850
rect 2090 -867 2094 -850
rect 2123 -867 2127 -850
rect 2187 -866 2191 -850
rect 2384 -861 2387 -540
rect 2453 -776 2462 -478
rect 2805 -515 2817 -440
rect 2487 -660 2764 -651
rect 2403 -785 2705 -776
rect 2403 -791 2679 -785
rect 2410 -803 2414 -791
rect 2454 -803 2458 -791
rect 2498 -803 2502 -791
rect 2542 -803 2546 -791
rect 2586 -803 2590 -791
rect 2630 -803 2634 -791
rect 2446 -818 2450 -807
rect 2490 -818 2494 -807
rect 2534 -818 2538 -807
rect 2578 -818 2582 -807
rect 2622 -818 2626 -807
rect 2446 -822 2626 -818
rect 2622 -856 2631 -822
rect 2666 -853 2670 -807
rect 2697 -831 2704 -785
rect 2802 -844 2817 -515
rect 2945 -800 2967 -662
rect 2965 -818 2967 -800
rect 3120 -844 3135 -454
rect 2408 -861 2417 -860
rect 2186 -867 2346 -866
rect 2056 -882 2346 -867
rect 2384 -869 2417 -861
rect 2458 -870 2462 -861
rect 2507 -871 2510 -862
rect 2548 -871 2553 -862
rect 2592 -872 2597 -864
rect 2588 -873 2597 -872
rect 2622 -865 2638 -856
rect 2666 -865 2678 -853
rect 2802 -856 3139 -844
rect 2186 -883 2346 -882
rect 2338 -925 2346 -883
rect 2622 -906 2626 -865
rect 2666 -906 2670 -865
rect 2450 -910 2454 -906
rect 2494 -910 2498 -906
rect 2538 -910 2542 -906
rect 2582 -910 2586 -906
rect 2410 -924 2414 -910
rect 2630 -924 2634 -910
rect 2407 -925 2683 -924
rect 1976 -949 2206 -938
rect 2338 -939 2683 -925
rect 1976 -992 1983 -949
rect 2042 -950 2206 -949
rect 2060 -983 2064 -950
rect 2094 -983 2098 -950
rect 2127 -983 2131 -950
rect 2159 -983 2163 -950
rect 2214 -964 2279 -958
rect 2214 -983 2218 -964
rect 2246 -983 2250 -964
rect 1975 -1145 1983 -992
rect 2059 -1027 2063 -1021
rect 1994 -1038 2036 -1035
rect 2083 -1072 2087 -987
rect 2117 -1022 2121 -987
rect 2150 -1011 2154 -987
rect 2182 -1011 2186 -987
rect 2274 -967 2279 -964
rect 2274 -973 2498 -967
rect 2191 -1011 2195 -987
rect 2223 -1011 2227 -987
rect 2150 -1015 2227 -1011
rect 2092 -1028 2099 -1022
rect 2117 -1028 2166 -1022
rect 2092 -1035 2095 -1028
rect 2117 -1072 2121 -1028
rect 2226 -1052 2230 -1047
rect 2274 -1057 2279 -973
rect 2491 -1027 2518 -1021
rect 2491 -1028 2522 -1027
rect 2182 -1061 2279 -1057
rect 2182 -1072 2186 -1061
rect 2246 -1072 2250 -1061
rect 2154 -1076 2159 -1072
rect 2218 -1076 2223 -1072
rect 2060 -1093 2064 -1076
rect 2094 -1093 2098 -1076
rect 2127 -1093 2131 -1076
rect 2191 -1093 2195 -1076
rect 2062 -1108 2210 -1093
rect 2539 -1141 2551 -974
rect 2802 -1127 2817 -856
rect 3120 -857 3135 -856
rect 2802 -1141 2816 -1127
rect 1975 -1156 2203 -1145
rect 1986 -1382 1997 -1156
rect 2039 -1157 2203 -1156
rect 2057 -1190 2061 -1157
rect 2091 -1190 2095 -1157
rect 2124 -1190 2128 -1157
rect 2156 -1190 2160 -1157
rect 2539 -1158 2816 -1141
rect 2211 -1171 2277 -1165
rect 2211 -1190 2215 -1171
rect 2243 -1190 2247 -1171
rect 2056 -1234 2060 -1228
rect 2012 -1245 2036 -1242
rect 2080 -1279 2084 -1194
rect 2114 -1229 2118 -1194
rect 2147 -1218 2151 -1194
rect 2179 -1218 2183 -1194
rect 2188 -1218 2192 -1194
rect 2220 -1218 2224 -1194
rect 2147 -1222 2224 -1218
rect 2271 -1210 2276 -1171
rect 2539 -1210 2551 -1158
rect 2802 -1159 2816 -1158
rect 2271 -1211 2551 -1210
rect 2271 -1219 2300 -1211
rect 2308 -1219 2551 -1211
rect 2089 -1235 2096 -1229
rect 2114 -1235 2163 -1229
rect 2090 -1239 2093 -1235
rect 2114 -1279 2118 -1235
rect 2223 -1259 2227 -1254
rect 2271 -1264 2276 -1219
rect 2179 -1268 2277 -1264
rect 2179 -1279 2183 -1268
rect 2243 -1279 2247 -1268
rect 2151 -1283 2156 -1279
rect 2215 -1283 2220 -1279
rect 2057 -1299 2061 -1283
rect 2060 -1300 2061 -1299
rect 2091 -1300 2095 -1283
rect 2124 -1300 2128 -1283
rect 2188 -1300 2192 -1283
rect 2060 -1306 2207 -1300
rect 3533 -1306 3538 -235
rect 2060 -1313 3538 -1306
rect 2714 -1345 3503 -1333
rect 2754 -1366 2755 -1361
rect 2764 -1366 2790 -1361
rect 2510 -1371 2516 -1368
rect 2640 -1371 2646 -1370
rect 2509 -1376 2646 -1371
rect 2510 -1382 2516 -1376
rect 2640 -1381 2646 -1376
rect 2891 -1372 2898 -1371
rect 3017 -1372 3024 -1371
rect 2891 -1375 3025 -1372
rect 2891 -1381 2898 -1375
rect 3017 -1381 3024 -1375
rect 1986 -1383 2083 -1382
rect 1986 -1384 2180 -1383
rect 2263 -1384 2535 -1382
rect 1986 -1390 2535 -1384
rect 2032 -1507 2040 -1390
rect 2084 -1399 2089 -1390
rect 2115 -1399 2120 -1390
rect 2148 -1399 2153 -1390
rect 2263 -1391 2535 -1390
rect 2635 -1388 2907 -1381
rect 3009 -1388 3285 -1381
rect 2263 -1397 2539 -1391
rect 2635 -1396 2911 -1388
rect 3009 -1391 3409 -1388
rect 3009 -1396 3285 -1391
rect 2103 -1428 2108 -1404
rect 2134 -1428 2139 -1404
rect 2103 -1434 2153 -1428
rect 2167 -1431 2172 -1404
rect 2270 -1409 2274 -1397
rect 2314 -1409 2318 -1397
rect 2358 -1409 2362 -1397
rect 2402 -1409 2406 -1397
rect 2446 -1409 2450 -1397
rect 2490 -1409 2494 -1397
rect 2642 -1408 2646 -1396
rect 2686 -1408 2690 -1396
rect 2730 -1408 2734 -1396
rect 2774 -1408 2778 -1396
rect 2818 -1408 2822 -1396
rect 2862 -1408 2866 -1396
rect 3016 -1408 3020 -1396
rect 3060 -1408 3064 -1396
rect 3104 -1408 3108 -1396
rect 3148 -1408 3152 -1396
rect 3192 -1408 3196 -1396
rect 3236 -1408 3240 -1396
rect 2306 -1424 2310 -1413
rect 2350 -1424 2354 -1413
rect 2394 -1424 2398 -1413
rect 2438 -1424 2442 -1413
rect 2482 -1424 2486 -1413
rect 2306 -1428 2486 -1424
rect 2167 -1432 2215 -1431
rect 2053 -1447 2090 -1442
rect 2053 -1489 2058 -1447
rect 2117 -1447 2121 -1442
rect 2134 -1457 2139 -1434
rect 2167 -1436 2216 -1432
rect 2167 -1457 2172 -1436
rect 2108 -1462 2115 -1457
rect 2084 -1466 2089 -1462
rect 2148 -1466 2153 -1462
rect 2085 -1473 2185 -1466
rect 2053 -1492 2205 -1489
rect 2086 -1507 2176 -1503
rect 2032 -1513 2176 -1507
rect 2104 -1525 2108 -1513
rect 2120 -1550 2122 -1546
rect 2152 -1547 2156 -1529
rect 2200 -1547 2205 -1492
rect 2152 -1553 2205 -1547
rect 2152 -1563 2156 -1553
rect -574 -1664 -552 -1574
rect 2104 -1592 2108 -1567
rect 2093 -1602 2170 -1592
rect 2110 -1664 2121 -1602
rect -574 -1676 2121 -1664
rect 2212 -1734 2216 -1436
rect 2482 -1462 2491 -1428
rect 2244 -1475 2277 -1466
rect 2313 -1468 2322 -1467
rect 2244 -1662 2248 -1475
rect 2317 -1476 2322 -1468
rect 2361 -1469 2370 -1468
rect 2366 -1477 2370 -1469
rect 2410 -1477 2413 -1468
rect 2452 -1479 2457 -1470
rect 2482 -1471 2498 -1462
rect 2526 -1470 2530 -1413
rect 2678 -1423 2682 -1412
rect 2722 -1423 2726 -1412
rect 2766 -1423 2770 -1412
rect 2810 -1423 2814 -1412
rect 2854 -1423 2858 -1412
rect 2678 -1427 2858 -1423
rect 2854 -1461 2863 -1427
rect 2898 -1457 2902 -1412
rect 3052 -1423 3056 -1412
rect 3096 -1423 3100 -1412
rect 3140 -1423 3144 -1412
rect 3184 -1423 3188 -1412
rect 3228 -1423 3232 -1412
rect 3052 -1427 3232 -1423
rect 2526 -1471 2538 -1470
rect 2482 -1512 2486 -1471
rect 2526 -1512 2530 -1471
rect 2310 -1516 2314 -1512
rect 2354 -1516 2358 -1512
rect 2398 -1516 2402 -1512
rect 2442 -1516 2446 -1512
rect 2607 -1475 2649 -1465
rect 2689 -1475 2694 -1466
rect 2270 -1526 2274 -1516
rect 2268 -1531 2274 -1526
rect 2490 -1530 2494 -1516
rect 2277 -1531 2543 -1530
rect 2268 -1536 2531 -1531
rect 2260 -1538 2531 -1536
rect 2259 -1544 2531 -1538
rect 2259 -1587 2267 -1544
rect 2277 -1545 2531 -1544
rect 2287 -1558 2577 -1549
rect 2607 -1556 2612 -1475
rect 2739 -1476 2742 -1467
rect 2781 -1476 2785 -1467
rect 2827 -1478 2829 -1469
rect 2854 -1470 2870 -1461
rect 2854 -1511 2858 -1470
rect 2898 -1471 2949 -1457
rect 3228 -1461 3237 -1427
rect 3272 -1458 3276 -1412
rect 3401 -1438 3408 -1391
rect 3464 -1438 3650 -1437
rect 3401 -1441 3650 -1438
rect 3464 -1445 3650 -1441
rect 3272 -1461 3284 -1458
rect 3476 -1460 3480 -1445
rect 3609 -1460 3613 -1445
rect 2898 -1511 2902 -1471
rect 2682 -1515 2686 -1511
rect 2726 -1515 2730 -1511
rect 2770 -1515 2774 -1511
rect 2814 -1515 2818 -1511
rect 2642 -1527 2646 -1515
rect 2862 -1529 2866 -1515
rect 2647 -1542 2908 -1529
rect 2639 -1544 2915 -1542
rect 2803 -1556 2806 -1555
rect 2287 -1559 2381 -1558
rect 2301 -1571 2305 -1559
rect 2349 -1592 2353 -1575
rect 2569 -1573 2576 -1558
rect 2607 -1562 2806 -1556
rect 2569 -1583 2775 -1573
rect 2788 -1583 2789 -1573
rect 2569 -1584 2576 -1583
rect 2259 -1640 2270 -1604
rect 2349 -1599 2404 -1592
rect 2709 -1595 2713 -1583
rect 2349 -1609 2353 -1599
rect 2301 -1638 2305 -1613
rect 2294 -1640 2366 -1638
rect 2259 -1647 2366 -1640
rect 2294 -1648 2380 -1647
rect 2397 -1662 2404 -1599
rect 2725 -1620 2727 -1616
rect 2757 -1617 2761 -1599
rect 2803 -1617 2806 -1562
rect 2757 -1623 2808 -1617
rect 2757 -1633 2761 -1623
rect 2709 -1662 2713 -1637
rect 2244 -1665 2404 -1662
rect 2397 -1666 2404 -1665
rect 2699 -1672 2775 -1662
rect 2939 -1698 2949 -1471
rect 2986 -1474 3023 -1469
rect 2986 -1560 2993 -1474
rect 3063 -1475 3068 -1466
rect 3113 -1476 3116 -1467
rect 3155 -1476 3159 -1467
rect 3185 -1468 3201 -1467
rect 3195 -1469 3201 -1468
rect 3195 -1478 3203 -1469
rect 3228 -1470 3244 -1461
rect 3272 -1470 3422 -1461
rect 3505 -1464 3510 -1460
rect 3539 -1464 3543 -1460
rect 3572 -1464 3576 -1460
rect 3228 -1511 3232 -1470
rect 3272 -1511 3276 -1470
rect 3410 -1490 3420 -1470
rect 3410 -1493 3582 -1490
rect 3480 -1505 3484 -1504
rect 3056 -1515 3060 -1511
rect 3100 -1515 3104 -1511
rect 3144 -1515 3148 -1511
rect 3188 -1515 3192 -1511
rect 3445 -1508 3484 -1505
rect 3445 -1510 3483 -1508
rect 3516 -1509 3519 -1505
rect 3579 -1504 3582 -1493
rect 3551 -1510 3552 -1506
rect 3016 -1529 3020 -1515
rect 3236 -1529 3240 -1515
rect 3013 -1530 3277 -1529
rect 3023 -1543 3277 -1530
rect 3023 -1544 3289 -1543
rect 2986 -1564 3242 -1560
rect 2986 -1566 3241 -1564
rect 3126 -1582 3216 -1572
rect 3136 -1594 3140 -1582
rect 3152 -1619 3154 -1615
rect 3184 -1616 3188 -1598
rect 3184 -1618 3192 -1616
rect 3238 -1618 3241 -1566
rect 3184 -1622 3241 -1618
rect 3184 -1632 3188 -1622
rect 3238 -1623 3241 -1622
rect 3136 -1661 3140 -1636
rect 3126 -1671 3203 -1661
rect 2939 -1713 3380 -1698
rect 3445 -1734 3451 -1510
rect 3601 -1505 3605 -1464
rect 3634 -1505 3638 -1464
rect 3584 -1511 3585 -1507
rect 3601 -1509 3617 -1505
rect 3634 -1509 3647 -1505
rect 3601 -1521 3605 -1509
rect 3501 -1525 3605 -1521
rect 3501 -1542 3505 -1525
rect 3535 -1542 3539 -1525
rect 3568 -1542 3572 -1525
rect 3601 -1542 3605 -1525
rect 3634 -1542 3638 -1509
rect 3476 -1551 3480 -1546
rect 3510 -1554 3514 -1546
rect 3543 -1554 3547 -1546
rect 3576 -1554 3580 -1546
rect 3609 -1554 3613 -1546
rect 3482 -1562 3659 -1554
rect 2212 -1740 3453 -1734
<< m2contact >>
rect 486 1997 495 2004
rect 519 2008 525 2013
rect 522 1983 527 1988
rect 604 2008 609 2013
rect 666 1994 675 2003
rect 708 1998 715 2003
rect 602 1970 607 1975
rect 659 1972 664 1977
rect 737 2008 743 2013
rect 822 2008 827 2013
rect 741 1980 746 1985
rect 882 1994 891 2005
rect 939 2000 946 2005
rect 820 1970 825 1975
rect 877 1972 882 1977
rect 970 2010 976 2015
rect 1055 2010 1060 2015
rect 1147 1996 1156 2006
rect 1199 2001 1206 2006
rect 975 1982 980 1987
rect 1053 1972 1058 1977
rect 1110 1974 1115 1979
rect 1230 2011 1236 2016
rect 1315 2011 1320 2016
rect 1420 1998 1432 2006
rect 1234 1984 1239 1989
rect 1313 1973 1318 1978
rect 1370 1975 1375 1980
rect 486 1954 495 1961
rect 443 1800 452 1805
rect -303 1752 -293 1765
rect 520 1800 525 1805
rect 564 1810 570 1815
rect 551 1799 556 1804
rect 633 1810 638 1815
rect 631 1772 636 1777
rect 688 1774 693 1779
rect 460 1606 474 1620
rect 701 1756 710 1764
rect 750 1795 755 1800
rect 781 1795 786 1800
rect 838 1806 846 1811
rect 941 1789 946 1794
rect 976 1793 984 1800
rect 742 1767 751 1775
rect 845 1768 854 1776
rect 888 1713 898 1720
rect 922 1761 931 1769
rect 945 1713 954 1720
rect 794 1656 800 1662
rect 527 1607 535 1614
rect 526 1543 534 1550
rect 558 1554 564 1559
rect 561 1543 566 1548
rect 643 1554 648 1559
rect 641 1516 646 1521
rect 698 1518 703 1523
rect 563 1472 568 1479
rect 1146 1797 1151 1802
rect 1190 1807 1196 1812
rect 1177 1796 1182 1801
rect 1259 1807 1264 1812
rect 1257 1769 1262 1774
rect 1314 1771 1319 1776
rect 1086 1603 1100 1617
rect 1327 1753 1336 1761
rect 1376 1792 1381 1797
rect 1407 1792 1412 1797
rect 1464 1803 1472 1808
rect 1567 1786 1572 1791
rect 1606 1790 1612 1795
rect 1368 1764 1377 1772
rect 1471 1765 1480 1773
rect 1514 1710 1524 1717
rect 1548 1758 1557 1766
rect 1571 1710 1580 1717
rect 1420 1653 1426 1659
rect 1153 1604 1161 1611
rect 1153 1538 1160 1547
rect 1184 1551 1190 1556
rect 1187 1540 1192 1545
rect 1269 1551 1274 1556
rect 1267 1513 1272 1518
rect 1324 1515 1329 1520
rect 1189 1469 1194 1476
rect 1746 1797 1751 1802
rect 1790 1807 1796 1812
rect 1777 1796 1782 1801
rect 1859 1807 1864 1812
rect 1857 1769 1862 1774
rect 1914 1771 1919 1776
rect 1686 1603 1700 1617
rect 1927 1753 1936 1761
rect 1976 1792 1981 1797
rect 2007 1792 2012 1797
rect 2064 1803 2072 1808
rect 2167 1786 2172 1791
rect 2206 1790 2211 1795
rect 1968 1764 1977 1772
rect 2071 1765 2080 1773
rect 2114 1710 2124 1717
rect 2148 1758 2157 1766
rect 2171 1710 2180 1717
rect 2020 1653 2026 1659
rect 1753 1604 1761 1611
rect 1753 1541 1761 1548
rect 1784 1551 1790 1556
rect 1787 1540 1792 1545
rect 1869 1551 1874 1556
rect 1867 1513 1872 1518
rect 1924 1515 1929 1520
rect 1789 1469 1794 1476
rect 2349 1800 2354 1805
rect 2393 1810 2399 1815
rect 2380 1799 2385 1804
rect 2462 1810 2467 1815
rect 2460 1772 2465 1777
rect 2517 1774 2522 1779
rect 2289 1606 2303 1620
rect 2530 1756 2539 1764
rect 2579 1795 2584 1800
rect 2610 1795 2615 1800
rect 2667 1806 2675 1811
rect 2770 1789 2775 1794
rect 2571 1767 2580 1775
rect 2674 1768 2683 1776
rect 2717 1713 2727 1720
rect 2751 1761 2760 1769
rect 2774 1713 2783 1720
rect 2623 1656 2629 1662
rect 2356 1607 2364 1614
rect 2356 1543 2363 1550
rect 2387 1554 2393 1559
rect 2390 1543 2395 1548
rect 2472 1554 2477 1559
rect 2470 1516 2475 1521
rect 2527 1518 2532 1523
rect 2392 1472 2397 1479
rect 159 1354 176 1374
rect 160 1191 176 1213
rect 475 1197 481 1204
rect -302 1140 -295 1150
rect -301 1097 -296 1102
rect -663 1057 -652 1066
rect -470 1057 -459 1066
rect -551 1008 -537 1017
rect -519 1008 -499 1018
rect -416 1028 -410 1033
rect -382 1028 -377 1033
rect -301 1039 -296 1045
rect -171 1075 -166 1080
rect -34 1078 -29 1083
rect -301 1029 -296 1034
rect -244 1029 -239 1034
rect -142 1029 -136 1035
rect -109 1030 -104 1035
rect -5 1028 1 1033
rect 28 1028 33 1033
rect 86 1039 95 1045
rect -416 907 -409 913
rect -381 908 -376 913
rect -313 919 -306 925
rect -270 908 -264 914
rect -236 909 -231 914
rect -170 920 -163 925
rect -142 912 -136 918
rect -107 912 -102 917
rect -36 922 -31 927
rect 3 911 9 916
rect 34 911 39 916
rect 102 922 108 928
rect -616 870 -602 884
rect -143 874 -135 880
rect 115 712 130 720
rect -122 654 -116 659
rect -969 424 -964 432
rect -1171 355 -1161 363
rect -1149 320 -1144 328
rect -961 384 -949 393
rect -1140 223 -1132 232
rect -1026 309 -1017 315
rect -967 321 -962 326
rect -958 283 -946 292
rect -511 565 -497 575
rect -779 338 -771 359
rect -289 630 -282 635
rect -394 582 -389 591
rect -363 585 -358 590
rect -152 627 -146 634
rect -260 585 -255 591
rect -225 586 -220 591
rect -13 632 -8 638
rect -124 586 -118 593
rect -90 587 -85 592
rect 541 1183 548 1188
rect 572 1193 578 1198
rect 657 1193 662 1198
rect 719 1179 728 1188
rect 761 1183 768 1188
rect 575 1161 581 1166
rect 655 1155 660 1160
rect 712 1157 717 1162
rect 790 1193 796 1198
rect 875 1193 880 1198
rect 793 1162 799 1167
rect 935 1179 944 1190
rect 992 1185 999 1190
rect 873 1155 878 1160
rect 930 1157 935 1162
rect 1023 1195 1029 1200
rect 1026 1170 1033 1175
rect 1108 1195 1113 1200
rect 1200 1181 1209 1191
rect 1252 1186 1259 1191
rect 1106 1157 1111 1162
rect 1163 1159 1168 1164
rect 1283 1196 1289 1201
rect 1368 1196 1373 1201
rect 1473 1183 1485 1191
rect 1286 1168 1293 1173
rect 1366 1158 1371 1163
rect 1423 1160 1428 1165
rect 573 985 578 990
rect 617 995 623 1000
rect 604 984 609 989
rect 686 995 691 1000
rect 684 957 689 962
rect 741 959 746 964
rect 513 791 527 805
rect 754 941 763 949
rect 803 980 808 985
rect 834 980 839 985
rect 891 991 899 996
rect 994 974 999 979
rect 1029 978 1037 985
rect 795 952 804 960
rect 898 953 907 961
rect 941 898 951 905
rect 975 946 984 954
rect 998 898 1007 905
rect 847 841 853 847
rect 580 792 588 799
rect 579 728 587 735
rect 611 739 617 744
rect 614 728 619 733
rect 696 739 701 744
rect 694 701 699 706
rect 751 703 756 708
rect 616 657 621 664
rect 1199 982 1204 987
rect 1243 992 1249 997
rect 1230 981 1235 986
rect 1312 992 1317 997
rect 1310 954 1315 959
rect 1367 956 1372 961
rect 1139 788 1153 802
rect 1380 938 1389 946
rect 1429 977 1434 982
rect 1460 977 1465 982
rect 1517 988 1525 993
rect 1620 971 1625 976
rect 1659 975 1665 980
rect 1421 949 1430 957
rect 1524 950 1533 958
rect 1567 895 1577 902
rect 1601 943 1610 951
rect 1624 895 1633 902
rect 1473 838 1479 844
rect 1206 789 1214 796
rect 1206 723 1213 732
rect 1237 736 1243 741
rect 1240 725 1245 730
rect 1322 736 1327 741
rect 1320 698 1325 703
rect 1377 700 1382 705
rect 1242 654 1247 661
rect 1799 982 1804 987
rect 1843 992 1849 997
rect 1830 981 1835 986
rect 1912 992 1917 997
rect 1910 954 1915 959
rect 1967 956 1972 961
rect 1739 788 1753 802
rect 1980 938 1989 946
rect 2029 977 2034 982
rect 2060 977 2065 982
rect 2117 988 2125 993
rect 2220 971 2225 976
rect 2259 975 2264 980
rect 2021 949 2030 957
rect 2124 950 2133 958
rect 2167 895 2177 902
rect 2201 943 2210 951
rect 2224 895 2233 902
rect 2073 838 2079 844
rect 1806 789 1814 796
rect 1806 726 1814 733
rect 1837 736 1843 741
rect 1840 725 1845 730
rect 1922 736 1927 741
rect 1920 698 1925 703
rect 1977 700 1982 705
rect 1842 654 1847 661
rect 2402 985 2407 990
rect 2446 995 2452 1000
rect 2433 984 2438 989
rect 2515 995 2520 1000
rect 2513 957 2518 962
rect 2570 959 2575 964
rect 2342 791 2356 805
rect 2583 941 2592 949
rect 2632 980 2637 985
rect 2663 980 2668 985
rect 2720 991 2728 996
rect 2823 974 2828 979
rect 2624 952 2633 960
rect 2727 953 2736 961
rect 2770 898 2780 905
rect 2804 946 2813 954
rect 2827 898 2836 905
rect 2676 841 2682 847
rect 2409 792 2417 799
rect 2409 728 2416 735
rect 2440 739 2446 744
rect 2443 728 2448 733
rect 2525 739 2530 744
rect 2523 701 2528 706
rect 2580 703 2585 708
rect 2445 657 2450 664
rect 12 584 18 591
rect 47 585 52 590
rect -399 465 -392 470
rect -362 465 -357 470
rect -303 476 -297 482
rect -250 466 -245 472
rect -217 466 -212 471
rect -155 476 -149 482
rect -122 468 -116 475
rect -88 469 -83 474
rect -25 480 -19 486
rect 20 467 25 473
rect 53 468 58 473
rect 115 479 121 485
rect -516 441 -503 447
rect -895 321 -890 326
rect -1104 223 -1096 231
rect -964 218 -959 225
rect -955 184 -943 193
rect -1013 173 -1007 179
rect -1174 134 -1163 143
rect -650 262 -639 272
rect -886 218 -881 225
rect -1055 103 -1043 108
rect -1013 102 -1008 109
rect -557 213 -548 220
rect -647 162 -634 177
rect -498 140 -484 148
rect -1062 75 -1051 84
rect -953 76 -941 85
rect -382 158 -376 167
rect -350 160 -345 165
rect -285 169 -275 178
rect -247 160 -241 166
rect -212 161 -207 166
rect -146 171 -136 180
rect -111 161 -106 167
rect -77 162 -72 167
rect -9 171 1 180
rect 27 160 32 166
rect 60 160 65 165
rect -383 40 -378 46
rect -349 40 -344 45
rect -283 50 -278 57
rect -236 40 -231 46
rect -204 41 -199 46
rect -140 51 -135 57
rect -108 43 -102 49
rect -75 44 -70 49
rect -8 55 -2 61
rect 35 43 40 49
rect 66 43 71 48
rect 132 54 138 61
rect -645 4 -636 16
rect -678 -234 -666 -207
rect -446 -310 -432 -300
rect -330 -292 -323 -283
rect -298 -290 -293 -285
rect -229 -280 -223 -272
rect -195 -288 -187 -280
rect -160 -289 -155 -284
rect -74 -278 -68 -271
rect -61 -289 -55 -283
rect -25 -288 -20 -283
rect 62 -277 69 -271
rect 82 -290 87 -285
rect 112 -290 117 -285
rect 175 -349 186 -342
rect -831 -413 -823 -403
rect -297 -410 -292 -405
rect -644 -438 -634 -424
rect -187 -409 -181 -403
rect -152 -409 -147 -404
rect -203 -423 -197 -417
rect -92 -399 -86 -393
rect -56 -406 -49 -400
rect -23 -406 -18 -401
rect 47 -395 53 -389
rect 87 -407 93 -401
rect 118 -407 123 -402
rect 179 -396 185 -391
rect -227 -444 -220 -439
rect -202 -444 -195 -439
rect -74 -444 -68 -438
rect -179 -518 -173 -511
rect -240 -575 -235 -569
rect 1767 -313 1775 -302
rect 2288 168 2296 176
rect 1790 2 1799 10
rect 2000 -1 2010 10
rect 2145 27 2155 35
rect 2053 -16 2059 -9
rect 2327 23 2337 31
rect 2596 -10 2602 -5
rect 2698 -13 2704 -7
rect 2880 -10 2886 -5
rect 2398 -19 2407 -13
rect 2921 -14 2931 -7
rect 2136 -58 2148 -51
rect 2883 -170 2890 -161
rect 3462 -182 3467 -175
rect 2494 -224 2504 -215
rect 2201 -251 2214 -240
rect 2250 -250 2262 -241
rect 2346 -251 2356 -242
rect 2393 -253 2403 -244
rect 2310 -283 2315 -278
rect 2479 -245 2486 -234
rect 2598 -248 2604 -242
rect 2642 -249 2649 -243
rect 2685 -253 2695 -241
rect 2774 -252 2783 -245
rect 2864 -245 2873 -234
rect 2735 -279 2742 -271
rect 2975 -249 2987 -240
rect 3020 -250 3031 -241
rect 3069 -251 3080 -240
rect 3115 -251 3123 -242
rect 3245 -244 3256 -234
rect 3157 -278 3163 -271
rect 2031 -329 2043 -322
rect 2137 -328 2149 -321
rect 2177 -313 2182 -298
rect 3492 -185 3498 -175
rect 3527 -184 3533 -178
rect 3519 -247 3529 -240
rect 393 -413 398 -404
rect 2197 -442 2210 -431
rect 432 -470 437 -465
rect -168 -583 -161 -576
rect -11 -574 -5 -568
rect 212 -584 220 -578
rect -64 -632 -59 -626
rect 157 -642 163 -637
rect 189 -641 195 -636
rect 1983 -477 1992 -466
rect 2050 -558 2058 -546
rect 1998 -572 2003 -567
rect 2032 -570 2037 -565
rect 2089 -570 2095 -565
rect 2084 -579 2092 -574
rect 2216 -579 2223 -574
rect 2029 -636 2050 -619
rect 2313 -664 2330 -645
rect 2050 -804 2055 -795
rect 1998 -816 2005 -810
rect 2039 -816 2046 -810
rect 2089 -816 2096 -811
rect 2083 -826 2091 -821
rect 2215 -826 2222 -821
rect 2362 -850 2369 -834
rect 2037 -882 2056 -866
rect 2474 -660 2487 -649
rect 2764 -662 2781 -645
rect 2697 -845 2705 -831
rect 3120 -454 3135 -434
rect 2944 -662 2967 -648
rect 2945 -818 2965 -800
rect 2446 -870 2458 -860
rect 2498 -872 2507 -861
rect 2539 -872 2548 -862
rect 2584 -872 2592 -858
rect 2054 -1031 2059 -1020
rect 1989 -1038 1994 -1032
rect 2036 -1040 2042 -1035
rect 2498 -973 2508 -959
rect 2092 -1040 2098 -1035
rect 2087 -1052 2095 -1047
rect 2219 -1052 2226 -1047
rect 2538 -974 2552 -956
rect 2479 -1028 2491 -1013
rect 2518 -1027 2525 -1013
rect 2043 -1109 2062 -1093
rect 2050 -1236 2056 -1226
rect 2007 -1245 2012 -1239
rect 2036 -1246 2042 -1239
rect 2300 -1219 2308 -1211
rect 2090 -1245 2096 -1239
rect 2084 -1259 2092 -1254
rect 2216 -1259 2223 -1254
rect 2041 -1313 2060 -1299
rect 2697 -1345 2714 -1326
rect 3503 -1345 3514 -1333
rect 2755 -1366 2764 -1359
rect 2790 -1366 2799 -1359
rect 2535 -1391 2543 -1382
rect 2907 -1388 2919 -1381
rect 2110 -1449 2117 -1442
rect 2078 -1473 2085 -1466
rect 2176 -1514 2187 -1503
rect 2115 -1551 2120 -1545
rect 2084 -1604 2093 -1592
rect 2170 -1606 2184 -1591
rect 2309 -1476 2317 -1468
rect 2359 -1477 2366 -1469
rect 2402 -1477 2410 -1468
rect 2444 -1479 2452 -1470
rect 2530 -1470 2544 -1459
rect 2680 -1475 2689 -1466
rect 2531 -1546 2545 -1531
rect 2276 -1560 2287 -1549
rect 2726 -1476 2739 -1467
rect 2767 -1477 2781 -1467
rect 2817 -1478 2827 -1469
rect 2633 -1542 2647 -1527
rect 2908 -1542 2922 -1527
rect 2254 -1604 2270 -1587
rect 2314 -1596 2319 -1591
rect 2775 -1583 2788 -1573
rect 2366 -1647 2380 -1632
rect 2719 -1623 2725 -1614
rect 2685 -1677 2699 -1662
rect 2775 -1673 2789 -1658
rect 3050 -1475 3063 -1466
rect 3100 -1476 3113 -1467
rect 3142 -1476 3155 -1467
rect 3183 -1478 3195 -1468
rect 3511 -1509 3516 -1502
rect 3546 -1510 3551 -1503
rect 3009 -1545 3023 -1530
rect 3277 -1543 3291 -1528
rect 3113 -1582 3126 -1572
rect 3146 -1620 3152 -1615
rect 3112 -1672 3126 -1657
rect 3203 -1674 3217 -1659
rect 3380 -1721 3410 -1688
rect 3579 -1511 3584 -1504
rect 3468 -1566 3482 -1551
<< metal2 >>
rect 1181 2078 1200 2079
rect 469 2072 1287 2078
rect 469 2016 475 2072
rect 422 2011 475 2016
rect 422 1961 428 2011
rect 469 2003 475 2011
rect 525 2008 604 2012
rect 469 1998 486 2003
rect 708 2003 712 2072
rect 743 2008 822 2012
rect 939 2005 943 2072
rect 976 2010 1055 2014
rect 1199 2006 1203 2072
rect 1236 2011 1315 2015
rect 891 1994 905 2005
rect 486 1983 522 1987
rect 607 1972 659 1975
rect 422 1954 486 1961
rect -302 1150 -295 1752
rect 422 1549 428 1954
rect 670 1874 675 1994
rect 707 1981 741 1984
rect 825 1972 877 1975
rect 901 1908 905 1994
rect 1432 1998 2455 2005
rect 940 1982 975 1985
rect 1058 1974 1110 1977
rect 1147 1932 1156 1996
rect 1198 1984 1234 1987
rect 1318 1975 1370 1978
rect 1147 1922 1785 1932
rect 901 1905 1233 1908
rect 551 1871 785 1874
rect 1229 1871 1233 1905
rect 1780 1871 1785 1922
rect 2443 1874 2450 1998
rect 2380 1871 2614 1874
rect 452 1800 520 1805
rect 520 1795 525 1800
rect 551 1804 555 1871
rect 570 1810 633 1814
rect 781 1800 785 1871
rect 1177 1868 1411 1871
rect 875 1835 946 1839
rect 875 1811 879 1835
rect 846 1806 879 1811
rect 669 1795 750 1799
rect 520 1792 673 1795
rect 941 1794 946 1835
rect 1119 1810 1125 1811
rect 1118 1802 1150 1803
rect 984 1793 1030 1800
rect 1118 1797 1146 1802
rect 636 1774 688 1777
rect 742 1762 751 1767
rect 710 1756 751 1762
rect 701 1755 751 1756
rect 846 1757 853 1768
rect 922 1757 931 1761
rect 846 1752 931 1757
rect 898 1713 945 1720
rect 474 1607 527 1612
rect 474 1606 533 1607
rect 564 1554 643 1558
rect 422 1543 526 1549
rect 528 1460 534 1543
rect 563 1479 566 1543
rect 646 1518 698 1521
rect 794 1460 800 1656
rect 1026 1547 1030 1793
rect 1146 1792 1151 1797
rect 1177 1801 1181 1868
rect 1196 1807 1259 1811
rect 1407 1797 1411 1868
rect 1777 1868 2011 1871
rect 1501 1832 1572 1836
rect 1501 1808 1505 1832
rect 1472 1803 1505 1808
rect 1295 1792 1376 1796
rect 1146 1789 1299 1792
rect 1567 1791 1572 1832
rect 1743 1797 1746 1802
rect 1606 1795 1648 1796
rect 1612 1790 1648 1795
rect 1262 1771 1314 1774
rect 1368 1759 1377 1764
rect 1336 1753 1377 1759
rect 1327 1752 1377 1753
rect 1472 1754 1479 1765
rect 1548 1754 1557 1758
rect 1472 1749 1557 1754
rect 1524 1710 1571 1717
rect 1100 1604 1153 1609
rect 1100 1603 1159 1604
rect 1190 1551 1269 1555
rect 1026 1539 1153 1547
rect 528 1456 800 1460
rect 1154 1457 1160 1538
rect 1189 1476 1192 1540
rect 1272 1515 1324 1518
rect 1420 1457 1426 1653
rect 1644 1547 1648 1790
rect 1746 1792 1751 1797
rect 1777 1801 1781 1868
rect 1796 1807 1859 1811
rect 2007 1797 2011 1868
rect 2101 1832 2172 1836
rect 2101 1808 2105 1832
rect 2072 1803 2105 1808
rect 1895 1792 1976 1796
rect 1746 1789 1899 1792
rect 2167 1791 2172 1832
rect 2262 1804 2349 1805
rect 2278 1800 2349 1804
rect 2278 1796 2354 1800
rect 2380 1804 2384 1871
rect 2399 1810 2462 1814
rect 2610 1800 2614 1871
rect 2704 1835 2775 1839
rect 2704 1811 2708 1835
rect 2675 1806 2708 1811
rect 2349 1795 2354 1796
rect 2498 1795 2579 1799
rect 2211 1790 2252 1794
rect 2349 1792 2502 1795
rect 2770 1794 2775 1835
rect 1862 1771 1914 1774
rect 1968 1759 1977 1764
rect 1936 1753 1977 1759
rect 1927 1752 1977 1753
rect 2072 1754 2079 1765
rect 2148 1754 2157 1758
rect 2072 1749 2157 1754
rect 2124 1710 2171 1717
rect 1700 1604 1753 1609
rect 1700 1603 1759 1604
rect 1790 1551 1869 1555
rect 1644 1541 1753 1547
rect 1154 1453 1426 1457
rect 1754 1457 1760 1541
rect 1789 1476 1792 1540
rect 1872 1515 1924 1518
rect 2020 1457 2026 1653
rect 2242 1550 2251 1790
rect 2465 1774 2517 1777
rect 2571 1762 2580 1767
rect 2539 1756 2580 1762
rect 2530 1755 2580 1756
rect 2675 1757 2682 1768
rect 2751 1757 2760 1761
rect 2675 1752 2760 1757
rect 2727 1713 2774 1720
rect 2303 1607 2356 1612
rect 2303 1606 2362 1607
rect 2393 1554 2472 1558
rect 2242 1545 2356 1550
rect 2242 1544 2251 1545
rect 1754 1453 2026 1457
rect 2357 1460 2363 1543
rect 2392 1479 2395 1543
rect 2475 1518 2527 1521
rect 2623 1460 2629 1656
rect 2357 1456 2629 1460
rect 241 1405 2262 1417
rect 160 1213 172 1354
rect -897 1132 -428 1140
rect -513 1109 131 1117
rect -513 1106 -42 1109
rect -18 1106 131 1109
rect -513 1068 -503 1106
rect -822 1058 -663 1065
rect -822 1057 -794 1058
rect -652 1058 -651 1065
rect -513 1027 -502 1068
rect -513 1018 -503 1027
rect -879 1017 -630 1018
rect -879 1008 -551 1017
rect -879 429 -874 1008
rect -568 1007 -540 1008
rect -514 1004 -503 1008
rect -513 959 -504 1004
rect -514 870 -503 959
rect -468 913 -461 1057
rect -426 1033 -421 1072
rect -382 1033 -377 1106
rect -301 1045 -296 1097
rect -244 1034 -239 1106
rect -171 1080 -166 1097
rect -109 1035 -104 1106
rect -34 1083 -29 1098
rect -426 1028 -416 1033
rect -410 1028 -409 1033
rect -159 1030 -142 1035
rect -468 907 -416 913
rect -381 870 -376 908
rect -313 879 -308 919
rect -301 879 -298 1029
rect -282 908 -270 914
rect -282 897 -278 908
rect -236 870 -231 909
rect -168 880 -163 920
rect -159 901 -154 1030
rect 28 1033 33 1106
rect 241 1046 251 1405
rect 522 1257 1340 1263
rect 522 1201 528 1257
rect 481 1197 528 1201
rect 475 1196 528 1197
rect 86 1045 253 1046
rect 95 1039 253 1045
rect 241 1038 251 1039
rect -24 1028 -5 1033
rect -142 880 -137 912
rect -107 870 -102 912
rect -36 882 -31 922
rect -24 915 -17 1028
rect -24 882 -16 915
rect -7 911 3 916
rect 9 911 10 916
rect -7 881 -1 911
rect 34 870 39 911
rect 103 880 107 922
rect -845 590 -644 599
rect -633 590 -630 599
rect -964 425 -874 429
rect -614 448 -603 870
rect -514 862 159 870
rect -299 685 -296 846
rect -277 847 -267 851
rect -271 691 -267 847
rect 310 836 434 848
rect -148 821 -133 826
rect -138 686 -133 821
rect -22 689 -17 803
rect -4 689 0 815
rect 310 720 317 836
rect 475 734 481 1196
rect 522 1188 528 1196
rect 578 1193 657 1197
rect 761 1188 765 1257
rect 796 1193 875 1197
rect 992 1190 996 1257
rect 1029 1195 1108 1199
rect 1252 1191 1256 1257
rect 1289 1196 1368 1200
rect 522 1183 541 1188
rect 944 1179 958 1190
rect 567 1161 575 1165
rect 660 1157 712 1160
rect 723 1059 728 1179
rect 799 1163 852 1164
rect 799 1162 845 1163
rect 794 1160 845 1162
rect 878 1157 930 1160
rect 954 1093 958 1179
rect 1485 1183 2508 1190
rect 1033 1170 1183 1173
rect 1111 1159 1163 1162
rect 1200 1117 1209 1181
rect 1293 1169 2482 1172
rect 1371 1160 1423 1163
rect 1200 1107 1838 1117
rect 954 1090 1286 1093
rect 604 1056 838 1059
rect 1282 1056 1286 1090
rect 1833 1056 1838 1107
rect 2496 1059 2503 1183
rect 3066 1107 3076 1167
rect 3114 1131 3118 1195
rect 3066 1095 3076 1097
rect 2433 1056 2667 1059
rect 542 990 578 994
rect 573 980 578 985
rect 604 989 608 1056
rect 623 995 686 999
rect 834 985 838 1056
rect 1230 1053 1464 1056
rect 928 1020 999 1024
rect 928 996 932 1020
rect 899 991 932 996
rect 722 980 803 984
rect 573 977 726 980
rect 994 979 999 1020
rect 1037 978 1083 985
rect 1194 982 1199 987
rect 689 959 741 962
rect 795 947 804 952
rect 763 941 804 947
rect 754 940 804 941
rect 899 942 906 953
rect 975 942 984 946
rect 899 937 984 942
rect 951 898 998 905
rect 527 792 580 797
rect 527 791 586 792
rect 617 739 696 743
rect 475 728 579 734
rect 130 713 319 720
rect 102 674 144 675
rect -494 666 150 674
rect -494 663 -299 666
rect -270 663 150 666
rect -494 575 -484 663
rect -406 589 -394 591
rect -411 583 -394 589
rect -389 583 -388 591
rect -363 590 -358 663
rect -289 635 -282 655
rect -225 591 -220 663
rect -152 634 -145 653
rect -146 627 -145 634
rect -128 654 -122 659
rect -137 592 -133 654
rect -127 605 -124 654
rect -137 591 -124 592
rect -293 588 -260 591
rect -146 587 -124 591
rect -497 565 -484 575
rect -614 447 -504 448
rect -614 441 -516 447
rect -614 392 -603 441
rect -495 427 -484 565
rect -144 491 -141 587
rect -90 592 -85 663
rect -13 658 -8 659
rect -13 638 -8 652
rect -16 584 12 590
rect 47 590 52 663
rect 102 662 144 663
rect 581 645 587 728
rect 616 664 619 728
rect 699 703 751 706
rect 847 645 853 841
rect 1079 732 1083 978
rect 1199 977 1204 982
rect 1230 986 1234 1053
rect 1249 992 1312 996
rect 1460 982 1464 1053
rect 1830 1053 2064 1056
rect 1554 1017 1625 1021
rect 1554 993 1558 1017
rect 1525 988 1558 993
rect 1348 977 1429 981
rect 1199 974 1352 977
rect 1620 976 1625 1017
rect 1796 982 1799 987
rect 1659 980 1701 981
rect 1665 975 1701 980
rect 1315 956 1367 959
rect 1421 944 1430 949
rect 1389 938 1430 944
rect 1380 937 1430 938
rect 1525 939 1532 950
rect 1601 939 1610 943
rect 1525 934 1610 939
rect 1577 895 1624 902
rect 1153 789 1206 794
rect 1153 788 1212 789
rect 1243 736 1322 740
rect 1079 724 1206 732
rect 581 641 853 645
rect 1207 642 1213 723
rect 1242 661 1245 725
rect 1325 700 1377 703
rect 1473 642 1479 838
rect 1697 732 1701 975
rect 1799 977 1804 982
rect 1830 986 1834 1053
rect 1849 992 1912 996
rect 2060 982 2064 1053
rect 2154 1017 2225 1021
rect 2154 993 2158 1017
rect 2125 988 2158 993
rect 1948 977 2029 981
rect 1799 974 1952 977
rect 2220 976 2225 1017
rect 2399 985 2402 990
rect 2402 980 2407 985
rect 2433 989 2437 1056
rect 2452 995 2515 999
rect 2663 985 2667 1056
rect 2757 1020 2828 1024
rect 2757 996 2761 1020
rect 2728 991 2761 996
rect 2551 980 2632 984
rect 2264 975 2305 979
rect 2402 977 2555 980
rect 2823 979 2828 1020
rect 1915 956 1967 959
rect 2021 944 2030 949
rect 1989 938 2030 944
rect 1980 937 2030 938
rect 2125 939 2132 950
rect 2201 939 2210 943
rect 2125 934 2210 939
rect 2177 895 2224 902
rect 1753 789 1806 794
rect 1753 788 1812 789
rect 1843 736 1922 740
rect 1697 726 1806 732
rect 1207 638 1479 642
rect 1807 642 1813 726
rect 1842 661 1845 725
rect 1925 700 1977 703
rect 2073 642 2079 838
rect 2295 735 2304 975
rect 2518 959 2570 962
rect 2624 947 2633 952
rect 2592 941 2633 947
rect 2583 940 2633 941
rect 2728 942 2735 953
rect 2804 942 2813 946
rect 2728 937 2813 942
rect 2780 898 2827 905
rect 2356 792 2409 797
rect 2356 791 2415 792
rect 2446 739 2525 743
rect 2295 730 2409 735
rect 2295 729 2304 730
rect 1807 638 2079 642
rect 2410 645 2416 728
rect 2445 664 2448 728
rect 2528 703 2580 706
rect 2676 645 2682 841
rect 2410 641 2682 645
rect -128 495 -124 498
rect -297 476 -291 482
rect -149 476 -146 482
rect -436 467 -399 470
rect -362 427 -357 465
rect -297 436 -292 476
rect -265 466 -250 472
rect -217 427 -212 466
rect -150 437 -146 476
rect -129 478 -124 495
rect -19 480 -14 486
rect -129 475 -121 478
rect -129 470 -122 475
rect -128 468 -122 470
rect -128 437 -125 468
rect -88 427 -83 469
rect -20 439 -14 480
rect 121 479 125 485
rect 6 468 20 473
rect 8 439 13 468
rect 53 427 58 468
rect 120 439 125 479
rect -495 419 178 427
rect -949 384 -603 392
rect -10 402 -9 408
rect 7 405 8 408
rect -903 383 -603 384
rect -1169 143 -1164 355
rect -1144 320 -1033 328
rect -962 321 -895 326
rect -1132 223 -1104 226
rect -1168 83 -1163 134
rect -1091 108 -1088 320
rect -1036 315 -1033 320
rect -1036 309 -1026 315
rect -873 292 -865 383
rect -946 284 -865 292
rect -959 218 -886 225
rect -1010 179 -1007 207
rect -873 192 -865 284
rect -780 338 -779 356
rect -780 246 -772 338
rect -647 272 -641 383
rect -285 262 -282 346
rect -268 265 -265 348
rect -138 262 -135 376
rect -125 263 -122 377
rect -10 269 -5 402
rect 7 262 13 405
rect -780 238 -548 246
rect -843 203 -707 210
rect -943 184 -865 192
rect -1013 109 -1010 173
rect -1091 103 -1055 108
rect -873 88 -865 184
rect -950 85 -864 88
rect -1168 76 -1062 83
rect -941 80 -864 85
rect -678 -207 -667 238
rect -557 220 -548 238
rect -481 238 163 249
rect -645 16 -637 162
rect -481 150 -471 238
rect -399 166 -395 195
rect -399 161 -382 166
rect -398 160 -382 161
rect -350 165 -345 238
rect -483 148 -471 150
rect -484 140 -471 148
rect -905 -269 -687 -260
rect -914 -270 -671 -269
rect -831 -403 -825 -333
rect -644 -424 -637 4
rect -482 2 -471 140
rect -283 113 -278 169
rect -267 125 -264 198
rect -258 167 -255 188
rect -258 166 -243 167
rect -212 166 -207 238
rect -258 160 -247 166
rect -267 124 -261 125
rect -267 121 -265 124
rect -145 122 -141 171
rect -77 167 -72 238
rect -128 161 -111 167
rect -8 131 -3 171
rect 10 160 27 165
rect 60 165 65 238
rect 1820 174 1826 177
rect 1820 170 2288 174
rect -8 127 1623 131
rect -145 117 1595 122
rect -283 108 1240 113
rect 1190 107 1240 108
rect -282 57 -279 58
rect -422 40 -383 45
rect -349 2 -344 40
rect -282 32 -279 50
rect -261 45 -236 46
rect -257 41 -236 45
rect -204 2 -199 41
rect -139 31 -136 51
rect -113 44 -108 49
rect -75 2 -70 44
rect -6 35 -3 55
rect 21 44 35 49
rect 66 2 71 43
rect 135 37 138 54
rect -482 -6 191 2
rect 12 -33 30 -29
rect -272 -109 -268 -75
rect -261 -126 -257 -51
rect -98 -54 -97 -47
rect -228 -187 -207 -184
rect -127 -187 -123 -55
rect -100 -176 -97 -54
rect -100 -180 -73 -176
rect -127 -192 -89 -187
rect -77 -189 -73 -180
rect 27 -187 30 -33
rect 69 -157 73 -16
rect 69 -165 233 -157
rect 27 -190 54 -187
rect -429 -212 215 -201
rect -429 -300 -419 -212
rect -396 -286 -391 -268
rect -396 -291 -330 -286
rect -298 -285 -293 -212
rect -223 -280 -222 -273
rect -432 -310 -419 -300
rect -644 -439 -637 -438
rect -430 -448 -419 -310
rect -297 -448 -292 -410
rect -226 -439 -222 -280
rect -210 -288 -195 -284
rect -160 -284 -155 -212
rect -218 -289 -188 -288
rect -83 -252 -77 -247
rect -83 -383 -79 -252
rect -69 -263 -66 -261
rect -69 -267 -57 -263
rect -188 -403 -184 -389
rect -188 -409 -187 -403
rect -202 -439 -198 -423
rect -152 -448 -147 -409
rect -86 -417 -83 -393
rect -73 -438 -69 -278
rect -61 -283 -57 -267
rect -25 -283 -20 -212
rect 69 -277 70 -271
rect -55 -389 -53 -384
rect -59 -400 -53 -389
rect -59 -406 -56 -400
rect -23 -448 -18 -406
rect 47 -415 50 -395
rect 65 -417 70 -277
rect 112 -285 117 -212
rect 79 -290 82 -285
rect 227 -328 233 -165
rect 76 -333 233 -328
rect 77 -402 82 -333
rect 186 -349 264 -344
rect 260 -366 264 -349
rect 180 -391 249 -390
rect 185 -396 249 -391
rect 77 -406 87 -402
rect 118 -448 123 -407
rect -430 -456 227 -448
rect 241 -466 249 -396
rect 260 -406 265 -366
rect 260 -411 393 -406
rect 260 -511 265 -411
rect 1232 -447 1239 107
rect 1573 -396 1585 117
rect 1609 -344 1621 127
rect 1793 10 1796 12
rect 1793 -13 1796 2
rect 1651 -311 1767 -305
rect 1609 -354 1675 -344
rect 1609 -355 1621 -354
rect 1573 -408 1700 -396
rect 1232 -454 1760 -447
rect 1234 -455 1760 -454
rect 424 -470 432 -465
rect 424 -472 427 -470
rect -173 -518 265 -511
rect -118 -519 265 -518
rect -11 -568 -6 -519
rect -248 -575 -240 -571
rect -248 -579 -245 -575
rect -248 -582 -168 -579
rect 212 -578 218 -519
rect -72 -632 -64 -627
rect 75 -642 157 -637
rect 187 -641 189 -637
rect 187 -645 190 -641
rect 1793 -1241 1796 -20
rect 1820 -35 1826 170
rect 1899 146 2593 155
rect 1820 -1035 1826 -50
rect 1899 -59 1905 146
rect 2883 109 2886 110
rect 1952 105 2889 109
rect 1899 -810 1905 -73
rect 1952 -78 1955 105
rect 1985 90 2254 92
rect 1983 79 2254 90
rect 1952 -569 1955 -92
rect 1983 -466 1990 79
rect 2249 75 2254 79
rect 2248 67 2254 75
rect 2248 31 2253 67
rect 2155 27 2327 31
rect 2010 -1 2058 3
rect 2053 -9 2058 -1
rect 2596 -5 2599 94
rect 2883 -5 2886 105
rect 2407 -19 2454 -14
rect 2399 -20 2454 -19
rect 2141 -306 2145 -58
rect 2449 -105 2454 -20
rect 2701 -72 2704 -13
rect 2931 -13 2963 -8
rect 2572 -77 2704 -72
rect 2250 -111 2454 -105
rect 2536 -106 2543 -104
rect 2200 -251 2201 -246
rect 2250 -241 2255 -111
rect 2395 -216 2399 -215
rect 2350 -220 2494 -216
rect 2350 -242 2354 -220
rect 2395 -244 2399 -220
rect 2200 -272 2207 -251
rect 2536 -240 2543 -119
rect 2486 -245 2543 -240
rect 2479 -246 2543 -245
rect 2572 -244 2575 -77
rect 2885 -220 2890 -170
rect 2774 -227 2890 -220
rect 2572 -248 2598 -244
rect 2295 -272 2324 -271
rect 2642 -272 2645 -249
rect 2200 -274 2645 -272
rect 2200 -275 2302 -274
rect 2320 -275 2645 -274
rect 2774 -245 2778 -227
rect 2959 -242 2963 -13
rect 3343 -164 3351 -119
rect 3343 -172 3466 -164
rect 3462 -175 3466 -172
rect 2873 -245 2911 -242
rect 2774 -253 2778 -252
rect 2141 -309 2177 -306
rect 2017 -322 2036 -319
rect 2141 -321 2145 -309
rect 2017 -329 2031 -322
rect 2017 -330 2036 -329
rect 1952 -572 1998 -569
rect 2017 -619 2023 -330
rect 2200 -431 2207 -275
rect 2312 -344 2315 -283
rect 2685 -352 2693 -253
rect 2680 -353 2693 -352
rect 2499 -357 2693 -353
rect 2736 -357 2742 -279
rect 2906 -355 2910 -245
rect 2959 -246 2975 -242
rect 2499 -493 2505 -357
rect 2906 -358 2988 -355
rect 2041 -557 2050 -550
rect 2037 -570 2089 -567
rect 2095 -570 2477 -565
rect 2092 -579 2216 -574
rect 2017 -633 2029 -619
rect 2019 -636 2029 -633
rect 2019 -646 2040 -636
rect 1899 -816 1998 -810
rect 1899 -817 2005 -816
rect 2020 -872 2027 -646
rect 2330 -660 2474 -653
rect 2330 -661 2487 -660
rect 2499 -736 2506 -493
rect 2781 -662 2944 -652
rect 3020 -652 3029 -250
rect 3256 -244 3338 -240
rect 3493 -243 3497 -185
rect 3527 -240 3530 -184
rect 3254 -245 3338 -244
rect 2967 -662 3030 -652
rect 3071 -736 3078 -251
rect 3120 -434 3123 -251
rect 3158 -376 3162 -278
rect 3331 -280 3337 -245
rect 3474 -246 3497 -243
rect 3331 -286 3429 -280
rect 3474 -351 3480 -246
rect 3529 -243 3530 -240
rect 3519 -279 3525 -247
rect 2499 -745 3085 -736
rect 2042 -804 2050 -798
rect 2046 -816 2089 -813
rect 2096 -816 2302 -811
rect 2091 -826 2215 -821
rect 2295 -839 2301 -816
rect 2020 -881 2037 -872
rect 1820 -1038 1989 -1035
rect 2020 -1095 2027 -881
rect 2294 -1020 2302 -839
rect 2369 -850 2453 -845
rect 2362 -851 2453 -850
rect 2446 -860 2453 -851
rect 2499 -861 2506 -745
rect 3071 -747 3078 -745
rect 2584 -845 2697 -838
rect 2584 -849 2705 -845
rect 2584 -858 2592 -849
rect 2498 -959 2505 -872
rect 2542 -956 2546 -872
rect 2497 -973 2498 -960
rect 2049 -1029 2054 -1023
rect 2294 -1024 2479 -1020
rect 2042 -1040 2092 -1036
rect 2324 -1037 2367 -1036
rect 2098 -1040 2367 -1037
rect 2095 -1052 2219 -1047
rect 2020 -1100 2032 -1095
rect 2020 -1109 2043 -1100
rect 1793 -1242 1979 -1241
rect 1793 -1244 2007 -1242
rect 1952 -1431 1955 -1244
rect 1970 -1245 2007 -1244
rect 2020 -1307 2027 -1109
rect 2039 -1234 2050 -1229
rect 2042 -1245 2090 -1242
rect 2042 -1246 2095 -1245
rect 2092 -1259 2216 -1254
rect 2020 -1313 2041 -1307
rect 2020 -1322 2031 -1313
rect 1952 -1435 2010 -1431
rect 2020 -1598 2027 -1322
rect 2081 -1434 2105 -1433
rect 2081 -1437 2107 -1434
rect 2103 -1442 2107 -1437
rect 2102 -1449 2110 -1442
rect 2304 -1465 2307 -1219
rect 2064 -1473 2078 -1468
rect 2304 -1468 2310 -1465
rect 2064 -1474 2081 -1473
rect 2064 -1598 2073 -1474
rect 2304 -1476 2309 -1468
rect 2361 -1469 2366 -1040
rect 2497 -1273 2503 -973
rect 2525 -1023 2608 -1022
rect 2525 -1027 2781 -1023
rect 2593 -1029 2781 -1027
rect 2497 -1275 2704 -1273
rect 2726 -1275 2731 -1274
rect 2497 -1278 2733 -1275
rect 2498 -1280 2733 -1278
rect 2699 -1281 2733 -1280
rect 2571 -1336 2578 -1334
rect 2571 -1342 2697 -1336
rect 2543 -1391 2550 -1385
rect 2546 -1446 2550 -1391
rect 2305 -1494 2311 -1476
rect 2402 -1449 2550 -1446
rect 2402 -1468 2408 -1449
rect 2445 -1470 2451 -1449
rect 2546 -1450 2550 -1449
rect 2571 -1464 2578 -1342
rect 2726 -1359 2731 -1281
rect 2726 -1365 2755 -1359
rect 2544 -1470 2579 -1464
rect 2726 -1467 2731 -1365
rect 2768 -1467 2781 -1029
rect 2949 -1250 2965 -818
rect 3183 -1197 3191 -586
rect 2949 -1257 2966 -1250
rect 2949 -1264 3148 -1257
rect 2951 -1266 3148 -1264
rect 2799 -1365 3113 -1359
rect 2915 -1446 2918 -1388
rect 2682 -1494 2685 -1475
rect 2817 -1450 2918 -1446
rect 2817 -1469 2820 -1450
rect 3049 -1475 3050 -1471
rect 3101 -1467 3109 -1365
rect 3142 -1467 3148 -1266
rect 3049 -1494 3056 -1475
rect 3183 -1468 3192 -1197
rect 3142 -1477 3148 -1476
rect 2305 -1498 3057 -1494
rect 3511 -1502 3514 -1345
rect 2229 -1505 2232 -1504
rect 2187 -1512 2232 -1505
rect 2107 -1550 2115 -1546
rect 2229 -1551 2232 -1512
rect 3544 -1510 3546 -1503
rect 2545 -1542 2633 -1532
rect 2922 -1537 3009 -1534
rect 3291 -1542 3462 -1536
rect 2229 -1558 2276 -1551
rect 3455 -1555 3461 -1542
rect 3455 -1563 3468 -1555
rect 2788 -1582 3113 -1575
rect 2020 -1603 2084 -1598
rect 2020 -1607 2027 -1603
rect 2184 -1602 2254 -1593
rect 2314 -1600 2317 -1596
rect 2309 -1603 2317 -1600
rect 2672 -1620 2719 -1616
rect 2725 -1620 2726 -1616
rect 3083 -1620 3146 -1615
rect 2380 -1645 2667 -1641
rect 2654 -1664 2660 -1645
rect 2654 -1672 2685 -1664
rect 2789 -1672 3112 -1665
rect 2789 -1673 3118 -1672
rect 3455 -1661 3461 -1563
rect 3217 -1668 3463 -1661
rect 3544 -1700 3550 -1510
rect 3410 -1711 3559 -1700
<< m3contact >>
rect 481 1983 486 1990
rect 699 1980 707 1985
rect 931 1981 940 1988
rect 1193 1984 1198 1992
rect 1118 1803 1125 1810
rect 1738 1797 1743 1802
rect 2262 1796 2278 1804
rect 2262 1405 2280 1417
rect -915 1126 -897 1145
rect -428 1130 -416 1140
rect -426 1072 -421 1079
rect -833 1057 -822 1065
rect -171 1097 -166 1102
rect -34 1098 -29 1103
rect -283 892 -277 897
rect -313 874 -308 879
rect -302 874 -297 879
rect -158 896 -151 901
rect -168 875 -163 880
rect -36 877 -30 882
rect -24 875 -16 882
rect -7 875 -1 881
rect 103 874 108 880
rect -855 590 -845 603
rect -644 590 -633 605
rect -302 846 -296 852
rect -282 845 -277 852
rect -155 821 -148 827
rect -299 679 -294 685
rect -271 684 -264 691
rect -6 815 3 821
rect -22 803 -14 810
rect 434 835 447 850
rect 3111 1195 3122 1210
rect 562 1161 567 1166
rect 845 1157 852 1163
rect 1183 1170 1189 1175
rect 2482 1168 2488 1174
rect 3059 1167 3077 1182
rect 3109 1119 3127 1131
rect 3059 1097 3079 1107
rect 534 990 542 996
rect 1189 982 1194 987
rect -138 681 -132 686
rect -26 681 -18 689
rect -4 682 4 689
rect -411 589 -406 598
rect -289 655 -282 660
rect -298 588 -293 593
rect -152 653 -145 659
rect -137 654 -132 659
rect -127 600 -121 605
rect -14 652 -8 658
rect -22 584 -16 591
rect 1791 982 1796 987
rect 2391 985 2399 990
rect -135 495 -128 502
rect -144 486 -139 491
rect -447 467 -436 475
rect -270 466 -265 472
rect -297 431 -292 436
rect -150 432 -145 437
rect -128 431 -123 437
rect 1 468 6 474
rect -20 433 -14 439
rect 8 431 13 439
rect 120 433 125 439
rect -9 402 -4 408
rect 8 405 14 411
rect -139 376 -134 383
rect -128 377 -121 384
rect -286 346 -280 352
rect -271 348 -263 357
rect -285 255 -280 262
rect -269 258 -262 265
rect -138 256 -132 262
rect -125 257 -116 263
rect -10 261 0 269
rect 7 256 13 262
rect -851 203 -843 210
rect -707 200 -695 212
rect -400 195 -394 204
rect -267 198 -261 203
rect -915 -269 -905 -255
rect -687 -269 -667 -258
rect -831 -333 -823 -323
rect -260 188 -255 194
rect -265 117 -260 124
rect -133 161 -128 167
rect 5 160 10 166
rect -427 40 -422 46
rect -262 40 -257 45
rect -282 27 -277 32
rect -119 44 -113 50
rect -139 26 -134 31
rect 16 44 21 50
rect -6 28 -1 35
rect 133 30 141 37
rect 68 -16 74 -11
rect 5 -33 12 -27
rect -262 -51 -256 -45
rect -272 -75 -266 -68
rect -272 -115 -266 -109
rect -127 -55 -120 -50
rect -103 -54 -98 -47
rect -261 -132 -255 -126
rect -234 -187 -228 -182
rect -207 -187 -201 -181
rect -89 -192 -83 -187
rect -77 -196 -71 -189
rect 54 -193 61 -184
rect -399 -268 -391 -259
rect -218 -288 -210 -280
rect -77 -252 -69 -247
rect -71 -261 -66 -256
rect -189 -389 -183 -383
rect -83 -389 -78 -383
rect -86 -424 -80 -417
rect -60 -389 -55 -383
rect 47 -421 53 -415
rect 74 -290 79 -285
rect 64 -424 74 -417
rect 241 -478 252 -466
rect 1792 -20 1800 -13
rect 1641 -316 1651 -303
rect 1675 -357 1691 -340
rect 1700 -411 1718 -394
rect 1760 -461 1778 -441
rect 422 -477 427 -472
rect -77 -632 -72 -626
rect 68 -642 75 -636
rect 187 -650 192 -645
rect 2593 146 2599 155
rect 1817 -50 1828 -35
rect 1896 -73 1907 -59
rect 2596 94 2601 99
rect 1946 -92 1957 -78
rect 2536 -119 2546 -106
rect 3341 -119 3352 -110
rect 2312 -350 2317 -344
rect 2736 -367 2745 -357
rect 2988 -358 2996 -351
rect 2033 -557 2041 -546
rect 2477 -571 2486 -558
rect 3429 -286 3440 -276
rect 3519 -286 3529 -279
rect 3474 -358 3480 -351
rect 3157 -381 3165 -376
rect 3168 -586 3212 -538
rect 2034 -804 2042 -792
rect 2039 -1029 2049 -1019
rect 2032 -1234 2039 -1226
rect 2010 -1436 2016 -1429
rect 2074 -1437 2081 -1428
rect 2101 -1552 2107 -1542
rect 2304 -1603 2309 -1598
rect 2665 -1620 2672 -1615
rect 3071 -1621 3083 -1609
<< metal3 >>
rect 1100 2407 1193 2408
rect -627 2401 1193 2407
rect -911 918 -904 1126
rect -912 601 -903 918
rect -913 591 -855 601
rect -912 353 -903 591
rect -913 320 -903 353
rect -831 471 -824 1057
rect -627 790 -621 2401
rect 1100 2400 1193 2401
rect 902 2367 935 2369
rect -579 2358 935 2367
rect -579 815 -571 2358
rect -560 2340 -553 2341
rect -560 2336 703 2340
rect -560 1026 -553 2336
rect -531 2312 496 2324
rect -561 995 -552 1026
rect -560 840 -553 995
rect -531 851 -522 2312
rect 489 2015 495 2312
rect 481 2012 495 2015
rect 481 1990 484 2012
rect 698 1985 703 2336
rect 931 1988 934 2358
rect 698 1980 699 1985
rect 1187 1984 1193 2400
rect -172 1907 -165 1908
rect -174 1905 732 1907
rect -174 1899 1127 1905
rect -172 1457 -165 1899
rect 1118 1810 1125 1899
rect -34 1737 1551 1738
rect 1740 1737 1743 1797
rect -34 1728 1743 1737
rect -34 1727 1551 1728
rect -172 1448 -164 1457
rect -171 1132 -164 1448
rect -426 1079 -421 1130
rect -171 1102 -166 1132
rect -34 1103 -27 1727
rect 2262 1417 2278 1796
rect 562 1273 565 1274
rect 3178 1273 3195 1277
rect 562 1269 3195 1273
rect 562 1166 565 1269
rect 3040 1267 3195 1269
rect 2468 1205 2561 1206
rect 2468 1202 3111 1205
rect 2468 1173 2472 1202
rect 3054 1200 3111 1202
rect 1189 1170 2472 1173
rect 2488 1168 3059 1172
rect 3055 1162 3160 1163
rect 852 1158 3160 1162
rect 3055 1157 3160 1158
rect -29 1098 -27 1103
rect 190 990 534 996
rect -313 851 -308 874
rect -300 852 -297 874
rect -282 852 -278 892
rect -531 845 -308 851
rect -167 840 -163 875
rect -560 835 -162 840
rect -560 834 -163 835
rect -155 827 -152 896
rect -36 815 -30 877
rect -579 806 -29 815
rect -22 810 -18 875
rect -6 821 -2 875
rect 103 790 107 874
rect -627 785 108 790
rect 190 775 196 990
rect 1189 929 1192 982
rect -289 770 196 775
rect 248 922 1192 929
rect -633 590 -411 596
rect -298 593 -295 679
rect -289 676 -281 770
rect 248 759 257 922
rect 1793 870 1796 982
rect 289 866 1799 870
rect 289 863 296 866
rect 1793 865 1796 866
rect -152 754 257 759
rect -152 753 256 754
rect -289 660 -282 676
rect -297 488 -294 588
rect -297 485 -283 488
rect -831 467 -447 471
rect -913 209 -904 320
rect -913 203 -851 209
rect -843 203 -842 209
rect -913 177 -904 203
rect -914 121 -904 177
rect -914 -255 -905 121
rect -914 -270 -905 -269
rect -831 46 -824 467
rect -296 341 -293 431
rect -286 352 -283 485
rect -270 472 -267 684
rect -152 682 -146 753
rect -14 744 -9 745
rect 290 744 296 863
rect 2395 851 2399 985
rect 434 850 2401 851
rect 447 847 2401 850
rect -14 739 297 744
rect -152 659 -147 682
rect -137 659 -134 681
rect -134 600 -127 604
rect -134 502 -131 600
rect -22 591 -19 681
rect -14 658 -9 739
rect 290 738 296 739
rect -22 497 -19 584
rect -22 494 -5 497
rect -269 357 -266 466
rect -149 371 -146 432
rect -139 383 -136 491
rect -126 384 -123 431
rect -19 395 -16 433
rect -9 408 -5 494
rect 1 474 4 682
rect 8 411 13 431
rect 121 409 124 433
rect 3074 412 3079 1097
rect 3056 409 3080 412
rect 121 406 3080 409
rect 3056 405 3080 406
rect 3119 396 3127 1119
rect 3056 395 3127 396
rect -20 390 3127 395
rect 3056 389 3121 390
rect 3148 371 3158 1157
rect -149 366 3158 371
rect -149 365 3157 366
rect 3178 343 3195 1267
rect 3047 341 3195 343
rect -296 333 3195 341
rect 3047 330 3195 333
rect -695 200 -400 202
rect -707 197 -400 200
rect -284 192 -281 255
rect -267 203 -263 258
rect -132 256 -130 262
rect -284 189 -260 192
rect -831 41 -427 46
rect -831 -323 -824 41
rect -282 -80 -279 27
rect -272 -68 -269 189
rect -133 167 -130 256
rect -260 117 -259 123
rect -262 45 -259 117
rect -133 69 -129 161
rect -133 66 -124 69
rect -261 -45 -258 40
rect -138 -62 -135 26
rect -127 -50 -124 66
rect -119 50 -116 257
rect -9 192 -5 261
rect 8 206 12 256
rect 8 201 20 206
rect -9 189 8 192
rect 5 166 8 189
rect -116 -41 -113 44
rect -4 -11 -1 28
rect -4 -39 0 -11
rect 5 -27 9 160
rect 17 50 20 201
rect 2596 99 2599 146
rect 17 -12 20 44
rect 17 -16 68 -12
rect 134 -14 138 30
rect 134 -20 1792 -14
rect 134 -21 1796 -20
rect 134 -23 138 -21
rect -116 -44 -99 -41
rect -103 -47 -99 -44
rect -5 -48 1817 -39
rect -138 -68 1896 -62
rect -282 -82 -63 -80
rect -282 -87 1946 -82
rect -282 -88 -279 -87
rect -84 -88 1946 -87
rect -233 -111 -213 -110
rect -266 -115 -213 -111
rect -261 -183 -257 -132
rect -261 -187 -234 -183
rect -667 -268 -399 -261
rect -667 -269 -392 -268
rect -219 -280 -214 -115
rect 2546 -119 3341 -110
rect -219 -287 -218 -280
rect -204 -386 -201 -187
rect -88 -257 -85 -192
rect -77 -247 -72 -196
rect 55 -249 58 -193
rect 55 -250 77 -249
rect 55 -252 78 -250
rect 67 -253 78 -252
rect -88 -261 -71 -257
rect 75 -285 78 -253
rect 3440 -286 3519 -280
rect -204 -389 -189 -386
rect -78 -388 -60 -384
rect -86 -549 -82 -424
rect -86 -554 -73 -549
rect -77 -626 -73 -554
rect 47 -647 50 -421
rect 68 -636 73 -424
rect 252 -477 422 -473
rect 47 -650 187 -647
rect 1643 -1227 1649 -316
rect 1674 -353 1675 -345
rect 1691 -346 1779 -345
rect 1691 -350 2312 -346
rect 1691 -351 2315 -350
rect 1691 -353 1779 -351
rect 1678 -1021 1688 -357
rect 1706 -358 1712 -357
rect 1706 -359 1773 -358
rect 1706 -363 2736 -359
rect 1706 -365 1773 -363
rect 1706 -382 1712 -365
rect 2996 -358 3474 -353
rect 1705 -394 1712 -382
rect 1766 -377 1774 -376
rect 1766 -380 3157 -377
rect 1705 -797 1712 -411
rect 1766 -441 1774 -380
rect 1766 -550 1774 -461
rect 2036 -539 2261 -535
rect 2036 -546 2040 -539
rect 1766 -555 2033 -550
rect 2256 -608 2261 -539
rect 3051 -562 3168 -560
rect 2486 -570 3168 -562
rect 2486 -571 3061 -570
rect 2256 -616 3085 -608
rect 2256 -617 2261 -616
rect 2393 -767 2671 -759
rect 2037 -781 2042 -780
rect 2393 -781 2400 -767
rect 2037 -787 2400 -781
rect 2037 -792 2042 -787
rect 2393 -788 2400 -787
rect 1705 -804 2034 -797
rect 2043 -1007 2046 -1006
rect 2043 -1011 2317 -1007
rect 2043 -1019 2046 -1011
rect 1678 -1022 1709 -1021
rect 1678 -1029 2039 -1022
rect 1678 -1030 2047 -1029
rect 1678 -1032 1709 -1030
rect 1643 -1234 2032 -1227
rect 1643 -1235 1840 -1234
rect 1695 -1544 1702 -1235
rect 2016 -1436 2074 -1433
rect 1695 -1550 2101 -1544
rect 1714 -1551 2101 -1550
rect 2304 -1589 2316 -1011
rect 2304 -1598 2309 -1589
rect 2665 -1615 2671 -767
rect 3073 -798 3084 -616
rect 3072 -828 3084 -798
rect 3072 -1609 3078 -828
<< labels >>
rlabel metal1 -1144 447 -1144 447 1 vdd
rlabel metal1 -1185 138 -1185 138 1 gnd
rlabel metal1 -1241 407 -1241 407 1 node_s0
rlabel metal1 -1244 187 -1244 187 1 node_s1
rlabel metal1 -261 912 -261 912 1 node_b1
rlabel metal1 -134 914 -134 914 1 node_b2
rlabel m2contact 8 913 8 913 1 node_b3
rlabel m2contact -2 1029 -2 1029 1 node_a3
rlabel metal1 701 1545 701 1545 1 node_sa0
rlabel metal1 1328 1544 1328 1544 1 node_sa1
rlabel metal1 1929 1541 1929 1541 1 node_sa2
rlabel metal1 2532 1545 2532 1545 1 node_sa3
rlabel metal1 2806 1795 2806 1795 1 node_sac
rlabel metal1 756 728 756 728 1 node_ss0
rlabel metal1 1381 726 1381 726 1 node_ss1
rlabel metal1 1982 727 1982 727 1 node_ss2
rlabel metal1 2585 730 2585 730 1 node_ss3
rlabel metal1 2859 980 2859 980 1 node_ssc
rlabel metal1 2669 -859 2669 -859 1 node_c2
rlabel metal1 3591 -180 3591 -180 1 node_c1
rlabel metal1 3642 -1507 3642 -1507 1 node_c3
rlabel metal1 -182 -562 -182 -562 1 node_r0
rlabel metal1 -6 -618 -6 -618 1 node_r1
rlabel metal1 490 -455 490 -455 1 node_r3
rlabel metal1 248 -628 248 -628 1 node_r2
rlabel m2contact -137 1032 -137 1032 1 node_a2
rlabel metal1 -272 1031 -272 1031 1 node_a1
rlabel metal1 -408 1031 -408 1031 1 node_a0
rlabel metal1 -408 910 -408 910 1 node_b0
<< end >>
