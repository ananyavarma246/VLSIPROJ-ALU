magic
tech scmos
timestamp 1700179625
<< nwell >>
rect -2907 512 -2832 534
rect -2637 507 -2562 529
rect -2382 513 -2307 535
rect -2114 513 -2039 535
rect -1555 358 -1377 393
rect -2761 301 -2486 342
rect -2379 301 -2104 342
rect -1997 301 -1722 342
rect -2939 239 -2839 269
rect -2923 -16 -2719 16
rect -2924 -263 -2720 -231
rect -2570 -319 -2295 -278
rect -2920 -489 -2716 -457
rect -2923 -696 -2719 -664
rect -2896 -906 -2796 -876
rect -2710 -925 -2435 -884
rect -2338 -924 -2063 -883
rect -1964 -924 -1689 -883
rect -1505 -969 -1327 -934
rect -2880 -1027 -2805 -1005
rect -2683 -1073 -2608 -1051
rect -2275 -1097 -2200 -1075
rect -1848 -1096 -1773 -1074
<< ntransistor >>
rect -2873 476 -2869 490
rect -2603 471 -2599 485
rect -2348 477 -2344 491
rect -2080 477 -2076 491
rect -1536 290 -1532 299
rect -1501 290 -1497 299
rect -1468 290 -1464 299
rect -1435 290 -1431 299
rect -1402 290 -1398 299
rect -2739 217 -2735 228
rect -2693 217 -2689 228
rect -2648 217 -2644 228
rect -2605 217 -2601 228
rect -2560 217 -2556 228
rect -2517 217 -2513 228
rect -2357 217 -2353 228
rect -2311 217 -2307 228
rect -2266 217 -2262 228
rect -2223 217 -2219 228
rect -2178 217 -2174 228
rect -2135 217 -2131 228
rect -1975 217 -1971 228
rect -1929 217 -1925 228
rect -1884 217 -1880 228
rect -1841 217 -1837 228
rect -1796 217 -1792 228
rect -1753 217 -1749 228
rect -2924 193 -2920 202
rect -2892 193 -2888 202
rect -2858 193 -2854 202
rect -2907 -91 -2904 -85
rect -2872 -91 -2869 -85
rect -2837 -91 -2834 -85
rect -2805 -91 -2802 -85
rect -2774 -91 -2771 -85
rect -2741 -91 -2738 -85
rect -2908 -338 -2905 -332
rect -2873 -338 -2870 -332
rect -2838 -338 -2835 -332
rect -2806 -338 -2803 -332
rect -2775 -338 -2772 -332
rect -2742 -338 -2739 -332
rect -2548 -403 -2544 -392
rect -2502 -403 -2498 -392
rect -2457 -403 -2453 -392
rect -2414 -403 -2410 -392
rect -2369 -403 -2365 -392
rect -2326 -403 -2322 -392
rect -2904 -564 -2901 -558
rect -2869 -564 -2866 -558
rect -2834 -564 -2831 -558
rect -2802 -564 -2799 -558
rect -2771 -564 -2768 -558
rect -2738 -564 -2735 -558
rect -2907 -771 -2904 -765
rect -2872 -771 -2869 -765
rect -2837 -771 -2834 -765
rect -2805 -771 -2802 -765
rect -2774 -771 -2771 -765
rect -2741 -771 -2738 -765
rect -2881 -952 -2877 -943
rect -2849 -952 -2845 -943
rect -2815 -952 -2811 -943
rect -2688 -1009 -2684 -998
rect -2642 -1009 -2638 -998
rect -2597 -1009 -2593 -998
rect -2554 -1009 -2550 -998
rect -2509 -1009 -2505 -998
rect -2466 -1009 -2462 -998
rect -2316 -1008 -2312 -997
rect -2270 -1008 -2266 -997
rect -2225 -1008 -2221 -997
rect -2182 -1008 -2178 -997
rect -2137 -1008 -2133 -997
rect -2094 -1008 -2090 -997
rect -1942 -1008 -1938 -997
rect -1896 -1008 -1892 -997
rect -1851 -1008 -1847 -997
rect -1808 -1008 -1804 -997
rect -1763 -1008 -1759 -997
rect -1720 -1008 -1716 -997
rect -1486 -1037 -1482 -1028
rect -1451 -1037 -1447 -1028
rect -1418 -1037 -1414 -1028
rect -1385 -1037 -1381 -1028
rect -1352 -1037 -1348 -1028
rect -2846 -1063 -2842 -1049
rect -2649 -1109 -2645 -1095
rect -2241 -1133 -2237 -1119
rect -1814 -1132 -1810 -1118
<< ptransistor >>
rect -2873 518 -2869 528
rect -2603 513 -2599 523
rect -2348 519 -2344 529
rect -2080 519 -2076 529
rect -1536 372 -1532 381
rect -1501 372 -1497 381
rect -1468 372 -1464 381
rect -1435 372 -1431 381
rect -1402 372 -1398 381
rect -2739 320 -2735 331
rect -2693 320 -2689 331
rect -2648 320 -2644 331
rect -2605 320 -2601 331
rect -2560 320 -2556 331
rect -2517 320 -2513 331
rect -2357 320 -2353 331
rect -2311 320 -2307 331
rect -2266 320 -2262 331
rect -2223 320 -2219 331
rect -2178 320 -2174 331
rect -2135 320 -2131 331
rect -1975 320 -1971 331
rect -1929 320 -1925 331
rect -1884 320 -1880 331
rect -1841 320 -1837 331
rect -1796 320 -1792 331
rect -1753 320 -1749 331
rect -2924 251 -2920 260
rect -2892 251 -2888 260
rect -2858 251 -2854 260
rect -2907 -2 -2904 4
rect -2872 -2 -2869 4
rect -2837 -2 -2834 4
rect -2805 -2 -2802 4
rect -2774 -2 -2771 4
rect -2741 -2 -2738 4
rect -2908 -249 -2905 -243
rect -2873 -249 -2870 -243
rect -2838 -249 -2835 -243
rect -2806 -249 -2803 -243
rect -2775 -249 -2772 -243
rect -2742 -249 -2739 -243
rect -2548 -300 -2544 -289
rect -2502 -300 -2498 -289
rect -2457 -300 -2453 -289
rect -2414 -300 -2410 -289
rect -2369 -300 -2365 -289
rect -2326 -300 -2322 -289
rect -2904 -475 -2901 -469
rect -2869 -475 -2866 -469
rect -2834 -475 -2831 -469
rect -2802 -475 -2799 -469
rect -2771 -475 -2768 -469
rect -2738 -475 -2735 -469
rect -2907 -682 -2904 -676
rect -2872 -682 -2869 -676
rect -2837 -682 -2834 -676
rect -2805 -682 -2802 -676
rect -2774 -682 -2771 -676
rect -2741 -682 -2738 -676
rect -2881 -894 -2877 -885
rect -2849 -894 -2845 -885
rect -2815 -894 -2811 -885
rect -2688 -906 -2684 -895
rect -2642 -906 -2638 -895
rect -2597 -906 -2593 -895
rect -2554 -906 -2550 -895
rect -2509 -906 -2505 -895
rect -2466 -906 -2462 -895
rect -2316 -905 -2312 -894
rect -2270 -905 -2266 -894
rect -2225 -905 -2221 -894
rect -2182 -905 -2178 -894
rect -2137 -905 -2133 -894
rect -2094 -905 -2090 -894
rect -1942 -905 -1938 -894
rect -1896 -905 -1892 -894
rect -1851 -905 -1847 -894
rect -1808 -905 -1804 -894
rect -1763 -905 -1759 -894
rect -1720 -905 -1716 -894
rect -1486 -955 -1482 -946
rect -1451 -955 -1447 -946
rect -1418 -955 -1414 -946
rect -1385 -955 -1381 -946
rect -1352 -955 -1348 -946
rect -2846 -1021 -2842 -1011
rect -2649 -1067 -2645 -1057
rect -2241 -1091 -2237 -1081
rect -1814 -1090 -1810 -1080
<< ndiffusion >>
rect -2893 486 -2873 490
rect -2897 476 -2873 486
rect -2869 486 -2849 490
rect -2869 476 -2845 486
rect -2368 487 -2348 491
rect -2623 481 -2603 485
rect -2627 471 -2603 481
rect -2599 481 -2579 485
rect -2599 471 -2575 481
rect -2372 477 -2348 487
rect -2344 487 -2324 491
rect -2344 477 -2320 487
rect -2100 487 -2080 491
rect -2104 477 -2080 487
rect -2076 487 -2056 491
rect -2076 477 -2052 487
rect -1544 295 -1536 299
rect -1548 290 -1536 295
rect -1532 295 -1523 299
rect -1532 290 -1519 295
rect -1510 295 -1501 299
rect -1514 290 -1501 295
rect -1497 295 -1489 299
rect -1497 290 -1485 295
rect -1477 295 -1468 299
rect -1481 290 -1468 295
rect -1464 295 -1456 299
rect -1464 290 -1452 295
rect -1444 295 -1435 299
rect -1448 290 -1435 295
rect -1431 295 -1423 299
rect -1431 290 -1419 295
rect -1411 295 -1402 299
rect -1415 290 -1402 295
rect -1398 295 -1390 299
rect -1398 290 -1386 295
rect -2751 224 -2739 228
rect -2755 217 -2739 224
rect -2735 224 -2719 228
rect -2735 217 -2715 224
rect -2707 224 -2693 228
rect -2711 217 -2693 224
rect -2689 224 -2675 228
rect -2689 217 -2671 224
rect -2663 224 -2648 228
rect -2667 217 -2648 224
rect -2644 224 -2631 228
rect -2644 217 -2627 224
rect -2619 224 -2605 228
rect -2623 217 -2605 224
rect -2601 224 -2587 228
rect -2601 217 -2583 224
rect -2575 224 -2560 228
rect -2579 217 -2560 224
rect -2556 224 -2543 228
rect -2556 217 -2539 224
rect -2531 224 -2517 228
rect -2535 217 -2517 224
rect -2513 224 -2499 228
rect -2513 217 -2495 224
rect -2369 224 -2357 228
rect -2373 217 -2357 224
rect -2353 224 -2337 228
rect -2353 217 -2333 224
rect -2325 224 -2311 228
rect -2329 217 -2311 224
rect -2307 224 -2293 228
rect -2307 217 -2289 224
rect -2281 224 -2266 228
rect -2285 217 -2266 224
rect -2262 224 -2249 228
rect -2262 217 -2245 224
rect -2237 224 -2223 228
rect -2241 217 -2223 224
rect -2219 224 -2205 228
rect -2219 217 -2201 224
rect -2193 224 -2178 228
rect -2197 217 -2178 224
rect -2174 224 -2161 228
rect -2174 217 -2157 224
rect -2149 224 -2135 228
rect -2153 217 -2135 224
rect -2131 224 -2117 228
rect -2131 217 -2113 224
rect -1987 224 -1975 228
rect -1991 217 -1975 224
rect -1971 224 -1955 228
rect -1971 217 -1951 224
rect -1943 224 -1929 228
rect -1947 217 -1929 224
rect -1925 224 -1911 228
rect -1925 217 -1907 224
rect -1899 224 -1884 228
rect -1903 217 -1884 224
rect -1880 224 -1867 228
rect -1880 217 -1863 224
rect -1855 224 -1841 228
rect -1859 217 -1841 224
rect -1837 224 -1823 228
rect -1837 217 -1819 224
rect -1811 224 -1796 228
rect -1815 217 -1796 224
rect -1792 224 -1779 228
rect -1792 217 -1775 224
rect -1767 224 -1753 228
rect -1771 217 -1753 224
rect -1749 224 -1735 228
rect -1749 217 -1731 224
rect -2928 197 -2924 202
rect -2933 193 -2924 197
rect -2920 197 -2914 202
rect -2920 193 -2909 197
rect -2897 197 -2892 202
rect -2902 193 -2892 197
rect -2888 197 -2883 202
rect -2888 193 -2878 197
rect -2864 197 -2858 202
rect -2869 193 -2858 197
rect -2854 197 -2850 202
rect -2854 193 -2845 197
rect -2913 -89 -2907 -85
rect -2917 -91 -2907 -89
rect -2904 -89 -2894 -85
rect -2904 -91 -2890 -89
rect -2879 -89 -2872 -85
rect -2883 -91 -2872 -89
rect -2869 -89 -2860 -85
rect -2869 -91 -2856 -89
rect -2846 -89 -2837 -85
rect -2850 -91 -2837 -89
rect -2834 -89 -2827 -85
rect -2834 -91 -2823 -89
rect -2814 -89 -2805 -85
rect -2818 -91 -2805 -89
rect -2802 -89 -2795 -85
rect -2802 -91 -2791 -89
rect -2782 -89 -2774 -85
rect -2786 -91 -2774 -89
rect -2771 -89 -2763 -85
rect -2771 -91 -2759 -89
rect -2750 -89 -2741 -85
rect -2754 -91 -2741 -89
rect -2738 -89 -2731 -85
rect -2738 -91 -2727 -89
rect -2914 -336 -2908 -332
rect -2918 -338 -2908 -336
rect -2905 -336 -2895 -332
rect -2905 -338 -2891 -336
rect -2880 -336 -2873 -332
rect -2884 -338 -2873 -336
rect -2870 -336 -2861 -332
rect -2870 -338 -2857 -336
rect -2847 -336 -2838 -332
rect -2851 -338 -2838 -336
rect -2835 -336 -2828 -332
rect -2835 -338 -2824 -336
rect -2815 -336 -2806 -332
rect -2819 -338 -2806 -336
rect -2803 -336 -2796 -332
rect -2803 -338 -2792 -336
rect -2783 -336 -2775 -332
rect -2787 -338 -2775 -336
rect -2772 -336 -2764 -332
rect -2772 -338 -2760 -336
rect -2751 -336 -2742 -332
rect -2755 -338 -2742 -336
rect -2739 -336 -2732 -332
rect -2739 -338 -2728 -336
rect -2560 -396 -2548 -392
rect -2564 -403 -2548 -396
rect -2544 -396 -2528 -392
rect -2544 -403 -2524 -396
rect -2516 -396 -2502 -392
rect -2520 -403 -2502 -396
rect -2498 -396 -2484 -392
rect -2498 -403 -2480 -396
rect -2472 -396 -2457 -392
rect -2476 -403 -2457 -396
rect -2453 -396 -2440 -392
rect -2453 -403 -2436 -396
rect -2428 -396 -2414 -392
rect -2432 -403 -2414 -396
rect -2410 -396 -2396 -392
rect -2410 -403 -2392 -396
rect -2384 -396 -2369 -392
rect -2388 -403 -2369 -396
rect -2365 -396 -2352 -392
rect -2365 -403 -2348 -396
rect -2340 -396 -2326 -392
rect -2344 -403 -2326 -396
rect -2322 -396 -2308 -392
rect -2322 -403 -2304 -396
rect -2910 -562 -2904 -558
rect -2914 -564 -2904 -562
rect -2901 -562 -2891 -558
rect -2901 -564 -2887 -562
rect -2876 -562 -2869 -558
rect -2880 -564 -2869 -562
rect -2866 -562 -2857 -558
rect -2866 -564 -2853 -562
rect -2843 -562 -2834 -558
rect -2847 -564 -2834 -562
rect -2831 -562 -2824 -558
rect -2831 -564 -2820 -562
rect -2811 -562 -2802 -558
rect -2815 -564 -2802 -562
rect -2799 -562 -2792 -558
rect -2799 -564 -2788 -562
rect -2779 -562 -2771 -558
rect -2783 -564 -2771 -562
rect -2768 -562 -2760 -558
rect -2768 -564 -2756 -562
rect -2747 -562 -2738 -558
rect -2751 -564 -2738 -562
rect -2735 -562 -2728 -558
rect -2735 -564 -2724 -562
rect -2913 -769 -2907 -765
rect -2917 -771 -2907 -769
rect -2904 -769 -2894 -765
rect -2904 -771 -2890 -769
rect -2879 -769 -2872 -765
rect -2883 -771 -2872 -769
rect -2869 -769 -2860 -765
rect -2869 -771 -2856 -769
rect -2846 -769 -2837 -765
rect -2850 -771 -2837 -769
rect -2834 -769 -2827 -765
rect -2834 -771 -2823 -769
rect -2814 -769 -2805 -765
rect -2818 -771 -2805 -769
rect -2802 -769 -2795 -765
rect -2802 -771 -2791 -769
rect -2782 -769 -2774 -765
rect -2786 -771 -2774 -769
rect -2771 -769 -2763 -765
rect -2771 -771 -2759 -769
rect -2750 -769 -2741 -765
rect -2754 -771 -2741 -769
rect -2738 -769 -2731 -765
rect -2738 -771 -2727 -769
rect -2885 -948 -2881 -943
rect -2890 -952 -2881 -948
rect -2877 -948 -2871 -943
rect -2877 -952 -2866 -948
rect -2854 -948 -2849 -943
rect -2859 -952 -2849 -948
rect -2845 -948 -2840 -943
rect -2845 -952 -2835 -948
rect -2821 -948 -2815 -943
rect -2826 -952 -2815 -948
rect -2811 -948 -2807 -943
rect -2811 -952 -2802 -948
rect -2700 -1002 -2688 -998
rect -2704 -1009 -2688 -1002
rect -2684 -1002 -2668 -998
rect -2684 -1009 -2664 -1002
rect -2656 -1002 -2642 -998
rect -2660 -1009 -2642 -1002
rect -2638 -1002 -2624 -998
rect -2638 -1009 -2620 -1002
rect -2612 -1002 -2597 -998
rect -2616 -1009 -2597 -1002
rect -2593 -1002 -2580 -998
rect -2593 -1009 -2576 -1002
rect -2568 -1002 -2554 -998
rect -2572 -1009 -2554 -1002
rect -2550 -1002 -2536 -998
rect -2550 -1009 -2532 -1002
rect -2524 -1002 -2509 -998
rect -2528 -1009 -2509 -1002
rect -2505 -1002 -2492 -998
rect -2505 -1009 -2488 -1002
rect -2480 -1002 -2466 -998
rect -2484 -1009 -2466 -1002
rect -2462 -1002 -2448 -998
rect -2462 -1009 -2444 -1002
rect -2328 -1001 -2316 -997
rect -2332 -1008 -2316 -1001
rect -2312 -1001 -2296 -997
rect -2312 -1008 -2292 -1001
rect -2284 -1001 -2270 -997
rect -2288 -1008 -2270 -1001
rect -2266 -1001 -2252 -997
rect -2266 -1008 -2248 -1001
rect -2240 -1001 -2225 -997
rect -2244 -1008 -2225 -1001
rect -2221 -1001 -2208 -997
rect -2221 -1008 -2204 -1001
rect -2196 -1001 -2182 -997
rect -2200 -1008 -2182 -1001
rect -2178 -1001 -2164 -997
rect -2178 -1008 -2160 -1001
rect -2152 -1001 -2137 -997
rect -2156 -1008 -2137 -1001
rect -2133 -1001 -2120 -997
rect -2133 -1008 -2116 -1001
rect -2108 -1001 -2094 -997
rect -2112 -1008 -2094 -1001
rect -2090 -1001 -2076 -997
rect -2090 -1008 -2072 -1001
rect -1954 -1001 -1942 -997
rect -1958 -1008 -1942 -1001
rect -1938 -1001 -1922 -997
rect -1938 -1008 -1918 -1001
rect -1910 -1001 -1896 -997
rect -1914 -1008 -1896 -1001
rect -1892 -1001 -1878 -997
rect -1892 -1008 -1874 -1001
rect -1866 -1001 -1851 -997
rect -1870 -1008 -1851 -1001
rect -1847 -1001 -1834 -997
rect -1847 -1008 -1830 -1001
rect -1822 -1001 -1808 -997
rect -1826 -1008 -1808 -1001
rect -1804 -1001 -1790 -997
rect -1804 -1008 -1786 -1001
rect -1778 -1001 -1763 -997
rect -1782 -1008 -1763 -1001
rect -1759 -1001 -1746 -997
rect -1759 -1008 -1742 -1001
rect -1734 -1001 -1720 -997
rect -1738 -1008 -1720 -1001
rect -1716 -1001 -1702 -997
rect -1716 -1008 -1698 -1001
rect -1494 -1032 -1486 -1028
rect -1498 -1037 -1486 -1032
rect -1482 -1032 -1473 -1028
rect -1482 -1037 -1469 -1032
rect -1460 -1032 -1451 -1028
rect -1464 -1037 -1451 -1032
rect -1447 -1032 -1439 -1028
rect -1447 -1037 -1435 -1032
rect -1427 -1032 -1418 -1028
rect -1431 -1037 -1418 -1032
rect -1414 -1032 -1406 -1028
rect -1414 -1037 -1402 -1032
rect -1394 -1032 -1385 -1028
rect -1398 -1037 -1385 -1032
rect -1381 -1032 -1373 -1028
rect -1381 -1037 -1369 -1032
rect -1361 -1032 -1352 -1028
rect -1365 -1037 -1352 -1032
rect -1348 -1032 -1340 -1028
rect -1348 -1037 -1336 -1032
rect -2866 -1053 -2846 -1049
rect -2870 -1063 -2846 -1053
rect -2842 -1053 -2822 -1049
rect -2842 -1063 -2818 -1053
rect -2669 -1099 -2649 -1095
rect -2673 -1109 -2649 -1099
rect -2645 -1099 -2625 -1095
rect -2645 -1109 -2621 -1099
rect -2261 -1123 -2241 -1119
rect -2265 -1133 -2241 -1123
rect -2237 -1123 -2217 -1119
rect -2237 -1133 -2213 -1123
rect -1834 -1122 -1814 -1118
rect -1838 -1132 -1814 -1122
rect -1810 -1122 -1790 -1118
rect -1810 -1132 -1786 -1122
<< pdiffusion >>
rect -2893 524 -2873 528
rect -2897 518 -2873 524
rect -2869 524 -2849 528
rect -2869 518 -2845 524
rect -2368 525 -2348 529
rect -2623 519 -2603 523
rect -2627 513 -2603 519
rect -2599 519 -2579 523
rect -2372 519 -2348 525
rect -2344 525 -2324 529
rect -2344 519 -2320 525
rect -2100 525 -2080 529
rect -2104 519 -2080 525
rect -2076 525 -2056 529
rect -2076 519 -2052 525
rect -2599 513 -2575 519
rect -1544 377 -1536 381
rect -1548 372 -1536 377
rect -1532 377 -1523 381
rect -1532 372 -1519 377
rect -1510 377 -1501 381
rect -1514 372 -1501 377
rect -1497 377 -1489 381
rect -1497 372 -1485 377
rect -1477 377 -1468 381
rect -1481 372 -1468 377
rect -1464 377 -1456 381
rect -1464 372 -1452 377
rect -1444 377 -1435 381
rect -1448 372 -1435 377
rect -1431 377 -1423 381
rect -1431 372 -1419 377
rect -1411 377 -1402 381
rect -1415 372 -1402 377
rect -1398 377 -1390 381
rect -1398 372 -1386 377
rect -2751 327 -2739 331
rect -2755 320 -2739 327
rect -2735 327 -2719 331
rect -2735 320 -2715 327
rect -2707 327 -2693 331
rect -2711 320 -2693 327
rect -2689 327 -2675 331
rect -2689 320 -2671 327
rect -2663 327 -2648 331
rect -2667 320 -2648 327
rect -2644 327 -2631 331
rect -2644 320 -2627 327
rect -2619 327 -2605 331
rect -2623 320 -2605 327
rect -2601 327 -2587 331
rect -2601 320 -2583 327
rect -2575 327 -2560 331
rect -2579 320 -2560 327
rect -2556 327 -2543 331
rect -2556 320 -2539 327
rect -2531 327 -2517 331
rect -2535 320 -2517 327
rect -2513 327 -2499 331
rect -2513 320 -2495 327
rect -2369 327 -2357 331
rect -2373 320 -2357 327
rect -2353 327 -2337 331
rect -2353 320 -2333 327
rect -2325 327 -2311 331
rect -2329 320 -2311 327
rect -2307 327 -2293 331
rect -2307 320 -2289 327
rect -2281 327 -2266 331
rect -2285 320 -2266 327
rect -2262 327 -2249 331
rect -2262 320 -2245 327
rect -2237 327 -2223 331
rect -2241 320 -2223 327
rect -2219 327 -2205 331
rect -2219 320 -2201 327
rect -2193 327 -2178 331
rect -2197 320 -2178 327
rect -2174 327 -2161 331
rect -2174 320 -2157 327
rect -2149 327 -2135 331
rect -2153 320 -2135 327
rect -2131 327 -2117 331
rect -2131 320 -2113 327
rect -1987 327 -1975 331
rect -1991 320 -1975 327
rect -1971 327 -1955 331
rect -1971 320 -1951 327
rect -1943 327 -1929 331
rect -1947 320 -1929 327
rect -1925 327 -1911 331
rect -1925 320 -1907 327
rect -1899 327 -1884 331
rect -1903 320 -1884 327
rect -1880 327 -1867 331
rect -1880 320 -1863 327
rect -1855 327 -1841 331
rect -1859 320 -1841 327
rect -1837 327 -1823 331
rect -1837 320 -1819 327
rect -1811 327 -1796 331
rect -1815 320 -1796 327
rect -1792 327 -1779 331
rect -1792 320 -1775 327
rect -1767 327 -1753 331
rect -1771 320 -1753 327
rect -1749 327 -1735 331
rect -1749 320 -1731 327
rect -2928 255 -2924 260
rect -2933 251 -2924 255
rect -2920 255 -2914 260
rect -2920 251 -2909 255
rect -2897 255 -2892 260
rect -2902 251 -2892 255
rect -2888 255 -2883 260
rect -2888 251 -2878 255
rect -2864 255 -2858 260
rect -2869 251 -2858 255
rect -2854 255 -2850 260
rect -2854 251 -2845 255
rect -2913 0 -2907 4
rect -2917 -2 -2907 0
rect -2904 0 -2894 4
rect -2904 -2 -2890 0
rect -2879 0 -2872 4
rect -2883 -2 -2872 0
rect -2869 0 -2860 4
rect -2869 -2 -2856 0
rect -2846 0 -2837 4
rect -2850 -2 -2837 0
rect -2834 0 -2827 4
rect -2834 -2 -2823 0
rect -2814 0 -2805 4
rect -2818 -2 -2805 0
rect -2802 0 -2795 4
rect -2802 -2 -2791 0
rect -2782 0 -2774 4
rect -2786 -2 -2774 0
rect -2771 0 -2763 4
rect -2771 -2 -2759 0
rect -2750 0 -2741 4
rect -2754 -2 -2741 0
rect -2738 0 -2731 4
rect -2738 -2 -2727 0
rect -2914 -247 -2908 -243
rect -2918 -249 -2908 -247
rect -2905 -247 -2895 -243
rect -2905 -249 -2891 -247
rect -2880 -247 -2873 -243
rect -2884 -249 -2873 -247
rect -2870 -247 -2861 -243
rect -2870 -249 -2857 -247
rect -2847 -247 -2838 -243
rect -2851 -249 -2838 -247
rect -2835 -247 -2828 -243
rect -2835 -249 -2824 -247
rect -2815 -247 -2806 -243
rect -2819 -249 -2806 -247
rect -2803 -247 -2796 -243
rect -2803 -249 -2792 -247
rect -2783 -247 -2775 -243
rect -2787 -249 -2775 -247
rect -2772 -247 -2764 -243
rect -2772 -249 -2760 -247
rect -2751 -247 -2742 -243
rect -2755 -249 -2742 -247
rect -2739 -247 -2732 -243
rect -2739 -249 -2728 -247
rect -2560 -293 -2548 -289
rect -2564 -300 -2548 -293
rect -2544 -293 -2528 -289
rect -2544 -300 -2524 -293
rect -2516 -293 -2502 -289
rect -2520 -300 -2502 -293
rect -2498 -293 -2484 -289
rect -2498 -300 -2480 -293
rect -2472 -293 -2457 -289
rect -2476 -300 -2457 -293
rect -2453 -293 -2440 -289
rect -2453 -300 -2436 -293
rect -2428 -293 -2414 -289
rect -2432 -300 -2414 -293
rect -2410 -293 -2396 -289
rect -2410 -300 -2392 -293
rect -2384 -293 -2369 -289
rect -2388 -300 -2369 -293
rect -2365 -293 -2352 -289
rect -2365 -300 -2348 -293
rect -2340 -293 -2326 -289
rect -2344 -300 -2326 -293
rect -2322 -293 -2308 -289
rect -2322 -300 -2304 -293
rect -2910 -473 -2904 -469
rect -2914 -475 -2904 -473
rect -2901 -473 -2891 -469
rect -2901 -475 -2887 -473
rect -2876 -473 -2869 -469
rect -2880 -475 -2869 -473
rect -2866 -473 -2857 -469
rect -2866 -475 -2853 -473
rect -2843 -473 -2834 -469
rect -2847 -475 -2834 -473
rect -2831 -473 -2824 -469
rect -2831 -475 -2820 -473
rect -2811 -473 -2802 -469
rect -2815 -475 -2802 -473
rect -2799 -473 -2792 -469
rect -2799 -475 -2788 -473
rect -2779 -473 -2771 -469
rect -2783 -475 -2771 -473
rect -2768 -473 -2760 -469
rect -2768 -475 -2756 -473
rect -2747 -473 -2738 -469
rect -2751 -475 -2738 -473
rect -2735 -473 -2728 -469
rect -2735 -475 -2724 -473
rect -2913 -680 -2907 -676
rect -2917 -682 -2907 -680
rect -2904 -680 -2894 -676
rect -2904 -682 -2890 -680
rect -2879 -680 -2872 -676
rect -2883 -682 -2872 -680
rect -2869 -680 -2860 -676
rect -2869 -682 -2856 -680
rect -2846 -680 -2837 -676
rect -2850 -682 -2837 -680
rect -2834 -680 -2827 -676
rect -2834 -682 -2823 -680
rect -2814 -680 -2805 -676
rect -2818 -682 -2805 -680
rect -2802 -680 -2795 -676
rect -2802 -682 -2791 -680
rect -2782 -680 -2774 -676
rect -2786 -682 -2774 -680
rect -2771 -680 -2763 -676
rect -2771 -682 -2759 -680
rect -2750 -680 -2741 -676
rect -2754 -682 -2741 -680
rect -2738 -680 -2731 -676
rect -2738 -682 -2727 -680
rect -2885 -890 -2881 -885
rect -2890 -894 -2881 -890
rect -2877 -890 -2871 -885
rect -2877 -894 -2866 -890
rect -2854 -890 -2849 -885
rect -2859 -894 -2849 -890
rect -2845 -890 -2840 -885
rect -2845 -894 -2835 -890
rect -2821 -890 -2815 -885
rect -2826 -894 -2815 -890
rect -2811 -890 -2807 -885
rect -2811 -894 -2802 -890
rect -2700 -899 -2688 -895
rect -2704 -906 -2688 -899
rect -2684 -899 -2668 -895
rect -2684 -906 -2664 -899
rect -2656 -899 -2642 -895
rect -2660 -906 -2642 -899
rect -2638 -899 -2624 -895
rect -2638 -906 -2620 -899
rect -2612 -899 -2597 -895
rect -2616 -906 -2597 -899
rect -2593 -899 -2580 -895
rect -2593 -906 -2576 -899
rect -2568 -899 -2554 -895
rect -2572 -906 -2554 -899
rect -2550 -899 -2536 -895
rect -2550 -906 -2532 -899
rect -2524 -899 -2509 -895
rect -2528 -906 -2509 -899
rect -2505 -899 -2492 -895
rect -2505 -906 -2488 -899
rect -2480 -899 -2466 -895
rect -2484 -906 -2466 -899
rect -2462 -899 -2448 -895
rect -2462 -906 -2444 -899
rect -2328 -898 -2316 -894
rect -2332 -905 -2316 -898
rect -2312 -898 -2296 -894
rect -2312 -905 -2292 -898
rect -2284 -898 -2270 -894
rect -2288 -905 -2270 -898
rect -2266 -898 -2252 -894
rect -2266 -905 -2248 -898
rect -2240 -898 -2225 -894
rect -2244 -905 -2225 -898
rect -2221 -898 -2208 -894
rect -2221 -905 -2204 -898
rect -2196 -898 -2182 -894
rect -2200 -905 -2182 -898
rect -2178 -898 -2164 -894
rect -2178 -905 -2160 -898
rect -2152 -898 -2137 -894
rect -2156 -905 -2137 -898
rect -2133 -898 -2120 -894
rect -2133 -905 -2116 -898
rect -2108 -898 -2094 -894
rect -2112 -905 -2094 -898
rect -2090 -898 -2076 -894
rect -2090 -905 -2072 -898
rect -1954 -898 -1942 -894
rect -1958 -905 -1942 -898
rect -1938 -898 -1922 -894
rect -1938 -905 -1918 -898
rect -1910 -898 -1896 -894
rect -1914 -905 -1896 -898
rect -1892 -898 -1878 -894
rect -1892 -905 -1874 -898
rect -1866 -898 -1851 -894
rect -1870 -905 -1851 -898
rect -1847 -898 -1834 -894
rect -1847 -905 -1830 -898
rect -1822 -898 -1808 -894
rect -1826 -905 -1808 -898
rect -1804 -898 -1790 -894
rect -1804 -905 -1786 -898
rect -1778 -898 -1763 -894
rect -1782 -905 -1763 -898
rect -1759 -898 -1746 -894
rect -1759 -905 -1742 -898
rect -1734 -898 -1720 -894
rect -1738 -905 -1720 -898
rect -1716 -898 -1702 -894
rect -1716 -905 -1698 -898
rect -1494 -950 -1486 -946
rect -1498 -955 -1486 -950
rect -1482 -950 -1473 -946
rect -1482 -955 -1469 -950
rect -1460 -950 -1451 -946
rect -1464 -955 -1451 -950
rect -1447 -950 -1439 -946
rect -1447 -955 -1435 -950
rect -1427 -950 -1418 -946
rect -1431 -955 -1418 -950
rect -1414 -950 -1406 -946
rect -1414 -955 -1402 -950
rect -1394 -950 -1385 -946
rect -1398 -955 -1385 -950
rect -1381 -950 -1373 -946
rect -1381 -955 -1369 -950
rect -1361 -950 -1352 -946
rect -1365 -955 -1352 -950
rect -1348 -950 -1340 -946
rect -1348 -955 -1336 -950
rect -2866 -1015 -2846 -1011
rect -2870 -1021 -2846 -1015
rect -2842 -1015 -2822 -1011
rect -2842 -1021 -2818 -1015
rect -2669 -1061 -2649 -1057
rect -2673 -1067 -2649 -1061
rect -2645 -1061 -2625 -1057
rect -2645 -1067 -2621 -1061
rect -2261 -1085 -2241 -1081
rect -2265 -1091 -2241 -1085
rect -2237 -1085 -2217 -1081
rect -2237 -1091 -2213 -1085
rect -1834 -1084 -1814 -1080
rect -1838 -1090 -1814 -1084
rect -1810 -1084 -1790 -1080
rect -1810 -1090 -1786 -1084
<< ndcontact >>
rect -2897 486 -2893 490
rect -2849 486 -2845 490
rect -2372 487 -2368 491
rect -2627 481 -2623 485
rect -2579 481 -2575 485
rect -2324 487 -2320 491
rect -2104 487 -2100 491
rect -2056 487 -2052 491
rect -1548 295 -1544 299
rect -1523 295 -1519 299
rect -1514 295 -1510 299
rect -1489 295 -1485 299
rect -1481 295 -1477 299
rect -1456 295 -1452 299
rect -1448 295 -1444 299
rect -1423 295 -1419 299
rect -1415 295 -1411 299
rect -1390 295 -1386 299
rect -2755 224 -2751 228
rect -2719 224 -2715 228
rect -2711 224 -2707 228
rect -2675 224 -2671 228
rect -2667 224 -2663 228
rect -2631 224 -2627 228
rect -2623 224 -2619 228
rect -2587 224 -2583 228
rect -2579 224 -2575 228
rect -2543 224 -2539 228
rect -2535 224 -2531 228
rect -2499 224 -2495 228
rect -2373 224 -2369 228
rect -2337 224 -2333 228
rect -2329 224 -2325 228
rect -2293 224 -2289 228
rect -2285 224 -2281 228
rect -2249 224 -2245 228
rect -2241 224 -2237 228
rect -2205 224 -2201 228
rect -2197 224 -2193 228
rect -2161 224 -2157 228
rect -2153 224 -2149 228
rect -2117 224 -2113 228
rect -1991 224 -1987 228
rect -1955 224 -1951 228
rect -1947 224 -1943 228
rect -1911 224 -1907 228
rect -1903 224 -1899 228
rect -1867 224 -1863 228
rect -1859 224 -1855 228
rect -1823 224 -1819 228
rect -1815 224 -1811 228
rect -1779 224 -1775 228
rect -1771 224 -1767 228
rect -1735 224 -1731 228
rect -2933 197 -2928 202
rect -2914 197 -2909 202
rect -2902 197 -2897 202
rect -2883 197 -2878 202
rect -2869 197 -2864 202
rect -2850 197 -2845 202
rect -2917 -89 -2913 -85
rect -2894 -89 -2890 -85
rect -2883 -89 -2879 -85
rect -2860 -89 -2856 -85
rect -2850 -89 -2846 -85
rect -2827 -89 -2823 -85
rect -2818 -89 -2814 -85
rect -2795 -89 -2791 -85
rect -2786 -89 -2782 -85
rect -2763 -89 -2759 -85
rect -2754 -89 -2750 -85
rect -2731 -89 -2727 -85
rect -2918 -336 -2914 -332
rect -2895 -336 -2891 -332
rect -2884 -336 -2880 -332
rect -2861 -336 -2857 -332
rect -2851 -336 -2847 -332
rect -2828 -336 -2824 -332
rect -2819 -336 -2815 -332
rect -2796 -336 -2792 -332
rect -2787 -336 -2783 -332
rect -2764 -336 -2760 -332
rect -2755 -336 -2751 -332
rect -2732 -336 -2728 -332
rect -2564 -396 -2560 -392
rect -2528 -396 -2524 -392
rect -2520 -396 -2516 -392
rect -2484 -396 -2480 -392
rect -2476 -396 -2472 -392
rect -2440 -396 -2436 -392
rect -2432 -396 -2428 -392
rect -2396 -396 -2392 -392
rect -2388 -396 -2384 -392
rect -2352 -396 -2348 -392
rect -2344 -396 -2340 -392
rect -2308 -396 -2304 -392
rect -2914 -562 -2910 -558
rect -2891 -562 -2887 -558
rect -2880 -562 -2876 -558
rect -2857 -562 -2853 -558
rect -2847 -562 -2843 -558
rect -2824 -562 -2820 -558
rect -2815 -562 -2811 -558
rect -2792 -562 -2788 -558
rect -2783 -562 -2779 -558
rect -2760 -562 -2756 -558
rect -2751 -562 -2747 -558
rect -2728 -562 -2724 -558
rect -2917 -769 -2913 -765
rect -2894 -769 -2890 -765
rect -2883 -769 -2879 -765
rect -2860 -769 -2856 -765
rect -2850 -769 -2846 -765
rect -2827 -769 -2823 -765
rect -2818 -769 -2814 -765
rect -2795 -769 -2791 -765
rect -2786 -769 -2782 -765
rect -2763 -769 -2759 -765
rect -2754 -769 -2750 -765
rect -2731 -769 -2727 -765
rect -2890 -948 -2885 -943
rect -2871 -948 -2866 -943
rect -2859 -948 -2854 -943
rect -2840 -948 -2835 -943
rect -2826 -948 -2821 -943
rect -2807 -948 -2802 -943
rect -2704 -1002 -2700 -998
rect -2668 -1002 -2664 -998
rect -2660 -1002 -2656 -998
rect -2624 -1002 -2620 -998
rect -2616 -1002 -2612 -998
rect -2580 -1002 -2576 -998
rect -2572 -1002 -2568 -998
rect -2536 -1002 -2532 -998
rect -2528 -1002 -2524 -998
rect -2492 -1002 -2488 -998
rect -2484 -1002 -2480 -998
rect -2448 -1002 -2444 -998
rect -2332 -1001 -2328 -997
rect -2296 -1001 -2292 -997
rect -2288 -1001 -2284 -997
rect -2252 -1001 -2248 -997
rect -2244 -1001 -2240 -997
rect -2208 -1001 -2204 -997
rect -2200 -1001 -2196 -997
rect -2164 -1001 -2160 -997
rect -2156 -1001 -2152 -997
rect -2120 -1001 -2116 -997
rect -2112 -1001 -2108 -997
rect -2076 -1001 -2072 -997
rect -1958 -1001 -1954 -997
rect -1922 -1001 -1918 -997
rect -1914 -1001 -1910 -997
rect -1878 -1001 -1874 -997
rect -1870 -1001 -1866 -997
rect -1834 -1001 -1830 -997
rect -1826 -1001 -1822 -997
rect -1790 -1001 -1786 -997
rect -1782 -1001 -1778 -997
rect -1746 -1001 -1742 -997
rect -1738 -1001 -1734 -997
rect -1702 -1001 -1698 -997
rect -1498 -1032 -1494 -1028
rect -1473 -1032 -1469 -1028
rect -1464 -1032 -1460 -1028
rect -1439 -1032 -1435 -1028
rect -1431 -1032 -1427 -1028
rect -1406 -1032 -1402 -1028
rect -1398 -1032 -1394 -1028
rect -1373 -1032 -1369 -1028
rect -1365 -1032 -1361 -1028
rect -1340 -1032 -1336 -1028
rect -2870 -1053 -2866 -1049
rect -2822 -1053 -2818 -1049
rect -2673 -1099 -2669 -1095
rect -2625 -1099 -2621 -1095
rect -2265 -1123 -2261 -1119
rect -2217 -1123 -2213 -1119
rect -1838 -1122 -1834 -1118
rect -1790 -1122 -1786 -1118
<< pdcontact >>
rect -2897 524 -2893 528
rect -2849 524 -2845 528
rect -2372 525 -2368 529
rect -2627 519 -2623 523
rect -2579 519 -2575 523
rect -2324 525 -2320 529
rect -2104 525 -2100 529
rect -2056 525 -2052 529
rect -1548 377 -1544 381
rect -1523 377 -1519 381
rect -1514 377 -1510 381
rect -1489 377 -1485 381
rect -1481 377 -1477 381
rect -1456 377 -1452 381
rect -1448 377 -1444 381
rect -1423 377 -1419 381
rect -1415 377 -1411 381
rect -1390 377 -1386 381
rect -2755 327 -2751 331
rect -2719 327 -2715 331
rect -2711 327 -2707 331
rect -2675 327 -2671 331
rect -2667 327 -2663 331
rect -2631 327 -2627 331
rect -2623 327 -2619 331
rect -2587 327 -2583 331
rect -2579 327 -2575 331
rect -2543 327 -2539 331
rect -2535 327 -2531 331
rect -2499 327 -2495 331
rect -2373 327 -2369 331
rect -2337 327 -2333 331
rect -2329 327 -2325 331
rect -2293 327 -2289 331
rect -2285 327 -2281 331
rect -2249 327 -2245 331
rect -2241 327 -2237 331
rect -2205 327 -2201 331
rect -2197 327 -2193 331
rect -2161 327 -2157 331
rect -2153 327 -2149 331
rect -2117 327 -2113 331
rect -1991 327 -1987 331
rect -1955 327 -1951 331
rect -1947 327 -1943 331
rect -1911 327 -1907 331
rect -1903 327 -1899 331
rect -1867 327 -1863 331
rect -1859 327 -1855 331
rect -1823 327 -1819 331
rect -1815 327 -1811 331
rect -1779 327 -1775 331
rect -1771 327 -1767 331
rect -1735 327 -1731 331
rect -2933 255 -2928 260
rect -2914 255 -2909 260
rect -2902 255 -2897 260
rect -2883 255 -2878 260
rect -2869 255 -2864 260
rect -2850 255 -2845 260
rect -2917 0 -2913 4
rect -2894 0 -2890 4
rect -2883 0 -2879 4
rect -2860 0 -2856 4
rect -2850 0 -2846 4
rect -2827 0 -2823 4
rect -2818 0 -2814 4
rect -2795 0 -2791 4
rect -2786 0 -2782 4
rect -2763 0 -2759 4
rect -2754 0 -2750 4
rect -2731 0 -2727 4
rect -2918 -247 -2914 -243
rect -2895 -247 -2891 -243
rect -2884 -247 -2880 -243
rect -2861 -247 -2857 -243
rect -2851 -247 -2847 -243
rect -2828 -247 -2824 -243
rect -2819 -247 -2815 -243
rect -2796 -247 -2792 -243
rect -2787 -247 -2783 -243
rect -2764 -247 -2760 -243
rect -2755 -247 -2751 -243
rect -2732 -247 -2728 -243
rect -2564 -293 -2560 -289
rect -2528 -293 -2524 -289
rect -2520 -293 -2516 -289
rect -2484 -293 -2480 -289
rect -2476 -293 -2472 -289
rect -2440 -293 -2436 -289
rect -2432 -293 -2428 -289
rect -2396 -293 -2392 -289
rect -2388 -293 -2384 -289
rect -2352 -293 -2348 -289
rect -2344 -293 -2340 -289
rect -2308 -293 -2304 -289
rect -2914 -473 -2910 -469
rect -2891 -473 -2887 -469
rect -2880 -473 -2876 -469
rect -2857 -473 -2853 -469
rect -2847 -473 -2843 -469
rect -2824 -473 -2820 -469
rect -2815 -473 -2811 -469
rect -2792 -473 -2788 -469
rect -2783 -473 -2779 -469
rect -2760 -473 -2756 -469
rect -2751 -473 -2747 -469
rect -2728 -473 -2724 -469
rect -2917 -680 -2913 -676
rect -2894 -680 -2890 -676
rect -2883 -680 -2879 -676
rect -2860 -680 -2856 -676
rect -2850 -680 -2846 -676
rect -2827 -680 -2823 -676
rect -2818 -680 -2814 -676
rect -2795 -680 -2791 -676
rect -2786 -680 -2782 -676
rect -2763 -680 -2759 -676
rect -2754 -680 -2750 -676
rect -2731 -680 -2727 -676
rect -2890 -890 -2885 -885
rect -2871 -890 -2866 -885
rect -2859 -890 -2854 -885
rect -2840 -890 -2835 -885
rect -2826 -890 -2821 -885
rect -2807 -890 -2802 -885
rect -2704 -899 -2700 -895
rect -2668 -899 -2664 -895
rect -2660 -899 -2656 -895
rect -2624 -899 -2620 -895
rect -2616 -899 -2612 -895
rect -2580 -899 -2576 -895
rect -2572 -899 -2568 -895
rect -2536 -899 -2532 -895
rect -2528 -899 -2524 -895
rect -2492 -899 -2488 -895
rect -2484 -899 -2480 -895
rect -2448 -899 -2444 -895
rect -2332 -898 -2328 -894
rect -2296 -898 -2292 -894
rect -2288 -898 -2284 -894
rect -2252 -898 -2248 -894
rect -2244 -898 -2240 -894
rect -2208 -898 -2204 -894
rect -2200 -898 -2196 -894
rect -2164 -898 -2160 -894
rect -2156 -898 -2152 -894
rect -2120 -898 -2116 -894
rect -2112 -898 -2108 -894
rect -2076 -898 -2072 -894
rect -1958 -898 -1954 -894
rect -1922 -898 -1918 -894
rect -1914 -898 -1910 -894
rect -1878 -898 -1874 -894
rect -1870 -898 -1866 -894
rect -1834 -898 -1830 -894
rect -1826 -898 -1822 -894
rect -1790 -898 -1786 -894
rect -1782 -898 -1778 -894
rect -1746 -898 -1742 -894
rect -1738 -898 -1734 -894
rect -1702 -898 -1698 -894
rect -1498 -950 -1494 -946
rect -1473 -950 -1469 -946
rect -1464 -950 -1460 -946
rect -1439 -950 -1435 -946
rect -1431 -950 -1427 -946
rect -1406 -950 -1402 -946
rect -1398 -950 -1394 -946
rect -1373 -950 -1369 -946
rect -1365 -950 -1361 -946
rect -1340 -950 -1336 -946
rect -2870 -1015 -2866 -1011
rect -2822 -1015 -2818 -1011
rect -2673 -1061 -2669 -1057
rect -2625 -1061 -2621 -1057
rect -2265 -1085 -2261 -1081
rect -2217 -1085 -2213 -1081
rect -1838 -1084 -1834 -1080
rect -1790 -1084 -1786 -1080
<< polysilicon >>
rect -2873 528 -2869 540
rect -2603 523 -2599 535
rect -2348 529 -2344 541
rect -2080 529 -2076 541
rect -2873 490 -2869 518
rect -2603 485 -2599 513
rect -2348 491 -2344 519
rect -2080 491 -2076 519
rect -2873 461 -2869 476
rect -2603 456 -2599 471
rect -2348 462 -2344 477
rect -2080 462 -2076 477
rect -1536 381 -1532 391
rect -1501 381 -1497 391
rect -1468 381 -1464 391
rect -1435 381 -1431 391
rect -1402 381 -1398 391
rect -2739 331 -2735 336
rect -2693 331 -2689 336
rect -2648 331 -2644 336
rect -2605 331 -2601 336
rect -2560 331 -2556 336
rect -2517 331 -2513 336
rect -2357 331 -2353 336
rect -2311 331 -2307 336
rect -2266 331 -2262 336
rect -2223 331 -2219 336
rect -2178 331 -2174 336
rect -2135 331 -2131 336
rect -1975 331 -1971 336
rect -1929 331 -1925 336
rect -1884 331 -1880 336
rect -1841 331 -1837 336
rect -1796 331 -1792 336
rect -1753 331 -1749 336
rect -2924 260 -2920 266
rect -2892 260 -2888 264
rect -2858 260 -2854 264
rect -2924 217 -2920 251
rect -2923 212 -2920 217
rect -2924 202 -2920 212
rect -2892 202 -2888 251
rect -2858 202 -2854 251
rect -2739 228 -2735 320
rect -2693 273 -2689 320
rect -2694 264 -2689 273
rect -2648 272 -2644 320
rect -2605 272 -2601 320
rect -2693 228 -2689 264
rect -2646 263 -2644 272
rect -2603 263 -2601 272
rect -2560 270 -2556 320
rect -2648 228 -2644 263
rect -2605 228 -2601 263
rect -2559 261 -2556 270
rect -2560 228 -2556 261
rect -2517 228 -2513 320
rect -2357 228 -2353 320
rect -2311 273 -2307 320
rect -2312 264 -2307 273
rect -2266 272 -2262 320
rect -2223 272 -2219 320
rect -2311 228 -2307 264
rect -2264 263 -2262 272
rect -2221 263 -2219 272
rect -2178 270 -2174 320
rect -2266 228 -2262 263
rect -2223 228 -2219 263
rect -2177 261 -2174 270
rect -2178 228 -2174 261
rect -2135 228 -2131 320
rect -1975 228 -1971 320
rect -1929 273 -1925 320
rect -1930 264 -1925 273
rect -1884 272 -1880 320
rect -1841 272 -1837 320
rect -1929 228 -1925 264
rect -1882 263 -1880 272
rect -1839 263 -1837 272
rect -1796 270 -1792 320
rect -1884 228 -1880 263
rect -1841 228 -1837 263
rect -1795 261 -1792 270
rect -1796 228 -1792 261
rect -1753 228 -1749 320
rect -1536 299 -1532 372
rect -1501 299 -1497 372
rect -1468 299 -1464 372
rect -1435 299 -1431 372
rect -1402 299 -1398 372
rect -1536 286 -1532 290
rect -1501 286 -1497 290
rect -1468 286 -1464 290
rect -1435 286 -1431 290
rect -1402 286 -1398 290
rect -2739 210 -2735 217
rect -2693 210 -2689 217
rect -2648 210 -2644 217
rect -2605 210 -2601 217
rect -2560 210 -2556 217
rect -2517 210 -2513 217
rect -2357 210 -2353 217
rect -2311 210 -2307 217
rect -2266 210 -2262 217
rect -2223 210 -2219 217
rect -2178 210 -2174 217
rect -2135 210 -2131 217
rect -1975 210 -1971 217
rect -1929 210 -1925 217
rect -1884 210 -1880 217
rect -1841 210 -1837 217
rect -1796 210 -1792 217
rect -1753 210 -1749 217
rect -2924 190 -2920 193
rect -2892 190 -2888 193
rect -2858 190 -2854 193
rect -2872 30 -2771 33
rect -2907 4 -2904 13
rect -2872 4 -2869 30
rect -2837 4 -2834 13
rect -2805 4 -2802 13
rect -2774 4 -2771 30
rect -2741 4 -2738 13
rect -2907 -85 -2904 -2
rect -2872 -85 -2869 -2
rect -2837 -85 -2834 -2
rect -2805 -85 -2802 -2
rect -2774 -85 -2771 -2
rect -2741 -85 -2738 -2
rect -2907 -102 -2904 -91
rect -2872 -99 -2869 -91
rect -2837 -102 -2834 -91
rect -2805 -99 -2802 -91
rect -2774 -99 -2771 -91
rect -2741 -99 -2738 -91
rect -2907 -104 -2834 -102
rect -2873 -217 -2772 -214
rect -2908 -243 -2905 -234
rect -2873 -243 -2870 -217
rect -2838 -243 -2835 -234
rect -2806 -243 -2803 -234
rect -2775 -243 -2772 -217
rect -2742 -243 -2739 -234
rect -2908 -332 -2905 -249
rect -2873 -332 -2870 -249
rect -2838 -332 -2835 -249
rect -2806 -332 -2803 -249
rect -2775 -332 -2772 -249
rect -2742 -332 -2739 -249
rect -2548 -289 -2544 -284
rect -2502 -289 -2498 -284
rect -2457 -289 -2453 -284
rect -2414 -289 -2410 -284
rect -2369 -289 -2365 -284
rect -2326 -289 -2322 -284
rect -2908 -349 -2905 -338
rect -2873 -346 -2870 -338
rect -2838 -349 -2835 -338
rect -2806 -346 -2803 -338
rect -2775 -346 -2772 -338
rect -2742 -346 -2739 -338
rect -2908 -351 -2835 -349
rect -2548 -392 -2544 -300
rect -2502 -347 -2498 -300
rect -2503 -356 -2498 -347
rect -2457 -348 -2453 -300
rect -2414 -348 -2410 -300
rect -2502 -392 -2498 -356
rect -2455 -357 -2453 -348
rect -2412 -357 -2410 -348
rect -2369 -350 -2365 -300
rect -2457 -392 -2453 -357
rect -2414 -392 -2410 -357
rect -2368 -359 -2365 -350
rect -2369 -392 -2365 -359
rect -2326 -392 -2322 -300
rect -2548 -410 -2544 -403
rect -2502 -410 -2498 -403
rect -2457 -410 -2453 -403
rect -2414 -410 -2410 -403
rect -2369 -410 -2365 -403
rect -2326 -410 -2322 -403
rect -2869 -443 -2768 -440
rect -2904 -469 -2901 -460
rect -2869 -469 -2866 -443
rect -2834 -469 -2831 -460
rect -2802 -469 -2799 -460
rect -2771 -469 -2768 -443
rect -2738 -469 -2735 -460
rect -2904 -558 -2901 -475
rect -2869 -558 -2866 -475
rect -2834 -558 -2831 -475
rect -2802 -558 -2799 -475
rect -2771 -558 -2768 -475
rect -2738 -558 -2735 -475
rect -2904 -575 -2901 -564
rect -2869 -572 -2866 -564
rect -2834 -575 -2831 -564
rect -2802 -572 -2799 -564
rect -2771 -572 -2768 -564
rect -2738 -572 -2735 -564
rect -2904 -577 -2831 -575
rect -2872 -650 -2771 -647
rect -2907 -676 -2904 -667
rect -2872 -676 -2869 -650
rect -2837 -676 -2834 -667
rect -2805 -676 -2802 -667
rect -2774 -676 -2771 -650
rect -2741 -676 -2738 -667
rect -2907 -765 -2904 -682
rect -2872 -765 -2869 -682
rect -2837 -765 -2834 -682
rect -2805 -765 -2802 -682
rect -2774 -765 -2771 -682
rect -2741 -765 -2738 -682
rect -2907 -782 -2904 -771
rect -2872 -779 -2869 -771
rect -2837 -782 -2834 -771
rect -2805 -779 -2802 -771
rect -2774 -779 -2771 -771
rect -2741 -779 -2738 -771
rect -2907 -784 -2834 -782
rect -2881 -885 -2877 -879
rect -2849 -885 -2845 -881
rect -2815 -885 -2811 -881
rect -2881 -928 -2877 -894
rect -2880 -933 -2877 -928
rect -2881 -943 -2877 -933
rect -2849 -943 -2845 -894
rect -2815 -943 -2811 -894
rect -2688 -895 -2684 -890
rect -2642 -895 -2638 -890
rect -2597 -895 -2593 -890
rect -2554 -895 -2550 -890
rect -2509 -895 -2505 -890
rect -2466 -895 -2462 -890
rect -2316 -894 -2312 -889
rect -2270 -894 -2266 -889
rect -2225 -894 -2221 -889
rect -2182 -894 -2178 -889
rect -2137 -894 -2133 -889
rect -2094 -894 -2090 -889
rect -1942 -894 -1938 -889
rect -1896 -894 -1892 -889
rect -1851 -894 -1847 -889
rect -1808 -894 -1804 -889
rect -1763 -894 -1759 -889
rect -1720 -894 -1716 -889
rect -2881 -955 -2877 -952
rect -2849 -955 -2845 -952
rect -2815 -955 -2811 -952
rect -2688 -998 -2684 -906
rect -2642 -953 -2638 -906
rect -2643 -962 -2638 -953
rect -2597 -954 -2593 -906
rect -2554 -954 -2550 -906
rect -2642 -998 -2638 -962
rect -2595 -963 -2593 -954
rect -2552 -963 -2550 -954
rect -2509 -956 -2505 -906
rect -2597 -998 -2593 -963
rect -2554 -998 -2550 -963
rect -2508 -965 -2505 -956
rect -2509 -998 -2505 -965
rect -2466 -998 -2462 -906
rect -2316 -997 -2312 -905
rect -2270 -952 -2266 -905
rect -2271 -961 -2266 -952
rect -2225 -953 -2221 -905
rect -2182 -953 -2178 -905
rect -2270 -997 -2266 -961
rect -2223 -962 -2221 -953
rect -2180 -962 -2178 -953
rect -2137 -955 -2133 -905
rect -2225 -997 -2221 -962
rect -2182 -997 -2178 -962
rect -2136 -964 -2133 -955
rect -2137 -997 -2133 -964
rect -2094 -997 -2090 -905
rect -1942 -997 -1938 -905
rect -1896 -952 -1892 -905
rect -1897 -961 -1892 -952
rect -1851 -953 -1847 -905
rect -1808 -953 -1804 -905
rect -1896 -997 -1892 -961
rect -1849 -962 -1847 -953
rect -1806 -962 -1804 -953
rect -1763 -955 -1759 -905
rect -1851 -997 -1847 -962
rect -1808 -997 -1804 -962
rect -1762 -964 -1759 -955
rect -1763 -997 -1759 -964
rect -1720 -997 -1716 -905
rect -1486 -946 -1482 -936
rect -1451 -946 -1447 -936
rect -1418 -946 -1414 -936
rect -1385 -946 -1381 -936
rect -1352 -946 -1348 -936
rect -2846 -1011 -2842 -999
rect -2688 -1016 -2684 -1009
rect -2642 -1016 -2638 -1009
rect -2597 -1016 -2593 -1009
rect -2554 -1016 -2550 -1009
rect -2509 -1016 -2505 -1009
rect -2466 -1016 -2462 -1009
rect -2316 -1015 -2312 -1008
rect -2270 -1015 -2266 -1008
rect -2225 -1015 -2221 -1008
rect -2182 -1015 -2178 -1008
rect -2137 -1015 -2133 -1008
rect -2094 -1015 -2090 -1008
rect -1942 -1015 -1938 -1008
rect -1896 -1015 -1892 -1008
rect -1851 -1015 -1847 -1008
rect -1808 -1015 -1804 -1008
rect -1763 -1015 -1759 -1008
rect -1720 -1015 -1716 -1008
rect -2846 -1049 -2842 -1021
rect -1486 -1028 -1482 -955
rect -1451 -1028 -1447 -955
rect -1418 -1028 -1414 -955
rect -1385 -1028 -1381 -955
rect -1352 -1028 -1348 -955
rect -1486 -1041 -1482 -1037
rect -1451 -1041 -1447 -1037
rect -1418 -1041 -1414 -1037
rect -1385 -1041 -1381 -1037
rect -1352 -1041 -1348 -1037
rect -2649 -1057 -2645 -1045
rect -2846 -1078 -2842 -1063
rect -2649 -1095 -2645 -1067
rect -2241 -1081 -2237 -1069
rect -1814 -1080 -1810 -1068
rect -2649 -1124 -2645 -1109
rect -2241 -1119 -2237 -1091
rect -1814 -1118 -1810 -1090
rect -2241 -1148 -2237 -1133
rect -1814 -1147 -1810 -1132
<< polycontact >>
rect -2879 503 -2873 507
rect -2609 498 -2603 502
rect -2354 504 -2348 508
rect -2086 504 -2080 508
rect -1540 333 -1536 337
rect -2748 265 -2739 274
rect -2927 212 -2923 217
rect -2896 212 -2892 217
rect -2864 225 -2858 231
rect -2703 264 -2694 273
rect -2655 263 -2646 272
rect -2612 263 -2603 272
rect -2568 261 -2559 270
rect -2527 269 -2517 278
rect -2366 265 -2357 274
rect -2321 264 -2312 273
rect -2273 263 -2264 272
rect -2230 263 -2221 272
rect -2186 261 -2177 270
rect -2145 269 -2135 278
rect -1984 265 -1975 274
rect -1939 264 -1930 273
rect -1891 263 -1882 272
rect -1848 263 -1839 272
rect -1804 261 -1795 270
rect -1763 269 -1753 278
rect -1505 332 -1501 336
rect -1472 331 -1468 335
rect -1439 330 -1435 334
rect -1407 332 -1402 336
rect -2914 -40 -2907 -34
rect -2878 -41 -2872 -35
rect -2811 -41 -2805 -35
rect -2747 -65 -2741 -60
rect -2915 -287 -2908 -281
rect -2879 -288 -2873 -282
rect -2812 -288 -2806 -282
rect -2748 -312 -2742 -307
rect -2557 -355 -2548 -346
rect -2512 -356 -2503 -347
rect -2464 -357 -2455 -348
rect -2421 -357 -2412 -348
rect -2377 -359 -2368 -350
rect -2336 -351 -2326 -342
rect -2911 -513 -2904 -507
rect -2875 -514 -2869 -508
rect -2808 -514 -2802 -508
rect -2744 -538 -2738 -533
rect -2914 -720 -2907 -714
rect -2878 -721 -2872 -715
rect -2811 -721 -2805 -715
rect -2747 -745 -2741 -740
rect -2884 -933 -2880 -928
rect -2853 -933 -2849 -928
rect -2821 -920 -2815 -914
rect -2697 -961 -2688 -952
rect -2652 -962 -2643 -953
rect -2604 -963 -2595 -954
rect -2561 -963 -2552 -954
rect -2517 -965 -2508 -956
rect -2476 -957 -2466 -948
rect -2325 -960 -2316 -951
rect -2280 -961 -2271 -952
rect -2232 -962 -2223 -953
rect -2189 -962 -2180 -953
rect -2145 -964 -2136 -955
rect -2104 -956 -2094 -947
rect -1951 -960 -1942 -951
rect -1906 -961 -1897 -952
rect -1858 -962 -1849 -953
rect -1815 -962 -1806 -953
rect -1771 -964 -1762 -955
rect -1730 -956 -1720 -947
rect -1490 -994 -1486 -990
rect -2852 -1036 -2846 -1032
rect -1455 -995 -1451 -991
rect -1422 -996 -1418 -992
rect -1389 -997 -1385 -993
rect -1357 -995 -1352 -991
rect -2655 -1082 -2649 -1078
rect -2247 -1106 -2241 -1102
rect -1820 -1105 -1814 -1101
<< metal1 >>
rect -2958 566 -2800 572
rect -2958 218 -2951 566
rect -2915 549 -2819 550
rect -2915 548 -2829 549
rect -2941 541 -2829 548
rect -2941 355 -2932 541
rect -2915 540 -2819 541
rect -2897 528 -2893 540
rect -2884 503 -2879 507
rect -2849 506 -2845 524
rect -2804 506 -2800 566
rect -2390 548 -2294 551
rect -2122 548 -2026 551
rect -2390 546 -2026 548
rect -2555 545 -2026 546
rect -2637 543 -2026 545
rect -2637 542 -2294 543
rect -2637 537 -2549 542
rect -2390 541 -2294 542
rect -2122 541 -2026 543
rect -2645 535 -2549 537
rect -2627 523 -2623 535
rect -2372 529 -2368 541
rect -2104 529 -2100 541
rect -2849 500 -2800 506
rect -2849 490 -2845 500
rect -2614 498 -2609 502
rect -2579 501 -2575 519
rect -2359 504 -2354 508
rect -2324 507 -2320 525
rect -2324 501 -2276 507
rect -2091 504 -2086 508
rect -2056 507 -2052 525
rect -2579 495 -2576 501
rect -2897 461 -2893 486
rect -2579 485 -2575 495
rect -2324 491 -2320 501
rect -2056 500 -2053 507
rect -2056 491 -2052 500
rect -2916 456 -2838 461
rect -2826 456 -2819 461
rect -2627 456 -2623 481
rect -2372 462 -2368 487
rect -2104 462 -2100 487
rect -2391 458 -2026 462
rect -2391 457 -2294 458
rect -2552 456 -2294 457
rect -2123 456 -2026 458
rect -2916 455 -2819 456
rect -2646 455 -2369 456
rect -2823 453 -2369 455
rect -2823 451 -2549 453
rect -2646 450 -2549 451
rect -1745 452 -1739 459
rect -1745 447 -1547 452
rect -1745 358 -1739 447
rect -1551 404 -1546 447
rect -1560 396 -1374 404
rect -1548 381 -1544 396
rect -1415 381 -1411 396
rect -1519 377 -1514 381
rect -1485 377 -1481 381
rect -1452 377 -1448 381
rect -2762 357 -2472 358
rect -2762 356 -2470 357
rect -2380 356 -1722 358
rect -2762 355 -1722 356
rect -2941 353 -1722 355
rect -2941 351 -2091 353
rect -2941 350 -2470 351
rect -2941 276 -2932 350
rect -2762 344 -2470 350
rect -2762 343 -2486 344
rect -2755 331 -2751 343
rect -2711 331 -2707 343
rect -2667 331 -2663 343
rect -2623 331 -2619 343
rect -2579 331 -2575 343
rect -2535 331 -2531 343
rect -2719 316 -2715 327
rect -2675 316 -2671 327
rect -2631 316 -2627 327
rect -2587 316 -2583 327
rect -2543 316 -2539 327
rect -2719 312 -2539 316
rect -2543 278 -2534 312
rect -2499 281 -2495 327
rect -2480 299 -2470 344
rect -2380 344 -2091 351
rect -2084 350 -1722 353
rect -2084 344 -2083 350
rect -2380 343 -2104 344
rect -1998 343 -1722 350
rect -2373 331 -2369 343
rect -2329 331 -2325 343
rect -2285 331 -2281 343
rect -2241 331 -2237 343
rect -2197 331 -2193 343
rect -2153 331 -2149 343
rect -1991 331 -1987 343
rect -1947 331 -1943 343
rect -1903 331 -1899 343
rect -1859 331 -1855 343
rect -1815 331 -1811 343
rect -1771 331 -1767 343
rect -1569 336 -1563 337
rect -1544 336 -1540 337
rect -1569 331 -1540 336
rect -1507 332 -1505 336
rect -2337 316 -2333 327
rect -2293 316 -2289 327
rect -2249 316 -2245 327
rect -2205 316 -2201 327
rect -2161 316 -2157 327
rect -2337 312 -2157 316
rect -2499 280 -2487 281
rect -2941 269 -2837 276
rect -2933 260 -2928 269
rect -2902 260 -2897 269
rect -2869 260 -2864 269
rect -2760 265 -2748 274
rect -2712 264 -2703 273
rect -2664 263 -2655 272
rect -2618 263 -2612 272
rect -2571 261 -2568 270
rect -2543 269 -2527 278
rect -2914 231 -2909 255
rect -2883 231 -2878 255
rect -2914 225 -2864 231
rect -2850 228 -2845 255
rect -2543 228 -2539 269
rect -2499 228 -2495 280
rect -2488 269 -2487 280
rect -2161 278 -2152 312
rect -2117 281 -2113 327
rect -1955 316 -1951 327
rect -1911 316 -1907 327
rect -1867 316 -1863 327
rect -1823 316 -1819 327
rect -1779 316 -1775 327
rect -1955 312 -1775 316
rect -2117 280 -2105 281
rect -2375 272 -2366 274
rect -2370 266 -2366 272
rect -2375 265 -2366 266
rect -2330 271 -2321 273
rect -2325 265 -2321 271
rect -2330 264 -2321 265
rect -2279 263 -2273 272
rect -2239 263 -2230 272
rect -2195 269 -2186 270
rect -2191 262 -2186 269
rect -2195 261 -2186 262
rect -2161 269 -2145 278
rect -2117 269 -2110 280
rect -1779 278 -1770 312
rect -1735 281 -1731 327
rect -1735 280 -1723 281
rect -2161 228 -2157 269
rect -2117 228 -2113 269
rect -1987 265 -1984 274
rect -1943 264 -1939 273
rect -1894 263 -1891 272
rect -1851 263 -1848 272
rect -1813 261 -1804 270
rect -1779 269 -1763 278
rect -1735 270 -1729 280
rect -1735 269 -1723 270
rect -1779 228 -1775 269
rect -1735 228 -1731 269
rect -2958 217 -2932 218
rect -2958 212 -2927 217
rect -2902 216 -2896 217
rect -2904 212 -2896 216
rect -2883 202 -2878 225
rect -2850 222 -2808 228
rect -2715 224 -2711 228
rect -2671 224 -2667 228
rect -2627 224 -2623 228
rect -2583 224 -2579 228
rect -2333 224 -2329 228
rect -2289 224 -2285 228
rect -2245 224 -2241 228
rect -2201 224 -2197 228
rect -1951 224 -1947 228
rect -1907 224 -1903 228
rect -1863 224 -1859 228
rect -1819 224 -1815 228
rect -2850 202 -2845 222
rect -2909 197 -2902 202
rect -2933 193 -2928 197
rect -2869 193 -2864 197
rect -2939 192 -2837 193
rect -2931 186 -2837 192
rect -2812 128 -2809 222
rect -2798 205 -2797 208
rect -2755 210 -2751 224
rect -2535 210 -2531 224
rect -2373 210 -2369 224
rect -2153 210 -2149 224
rect -1991 210 -1987 224
rect -1771 210 -1767 224
rect -2758 208 -2482 210
rect -2792 205 -2482 208
rect -2758 199 -2482 205
rect -2376 201 -2100 210
rect -1994 201 -1718 210
rect -2376 199 -1718 201
rect -2758 197 -1718 199
rect -2758 195 -2100 197
rect -1994 195 -1718 197
rect -1569 128 -1563 331
rect -1423 336 -1419 377
rect -1390 336 -1386 377
rect -1476 335 -1473 336
rect -1476 331 -1472 335
rect -1476 330 -1473 331
rect -1441 330 -1439 334
rect -1423 332 -1407 336
rect -1390 332 -1377 336
rect -1423 320 -1419 332
rect -1523 316 -1419 320
rect -1523 299 -1519 316
rect -1489 299 -1485 316
rect -1456 299 -1452 316
rect -1423 299 -1419 316
rect -1390 299 -1386 332
rect -1548 287 -1544 295
rect -1514 287 -1510 295
rect -1481 287 -1477 295
rect -1448 287 -1444 295
rect -1415 287 -1411 295
rect -1551 279 -1367 287
rect -2812 127 -2782 128
rect -2769 127 -1563 128
rect -2812 123 -1563 127
rect -2812 122 -2782 123
rect -2769 122 -1563 123
rect -2687 79 -2155 80
rect -2764 74 -2155 79
rect -2935 48 -2771 49
rect -2998 -198 -2991 48
rect -2982 37 -2512 48
rect -2917 4 -2913 37
rect -2883 4 -2879 37
rect -2850 4 -2846 37
rect -2818 4 -2814 37
rect -2795 36 -2512 37
rect -2763 23 -2699 29
rect -2763 4 -2759 23
rect -2731 4 -2727 23
rect -2922 -40 -2914 -34
rect -2894 -85 -2890 0
rect -2860 -35 -2856 0
rect -2827 -24 -2823 0
rect -2795 -24 -2791 0
rect -2786 -24 -2782 0
rect -2754 -24 -2750 0
rect -2703 -21 -2699 23
rect -2827 -28 -2750 -24
rect -2704 -26 -2587 -21
rect -2885 -41 -2878 -35
rect -2860 -41 -2811 -35
rect -2860 -85 -2856 -41
rect -2751 -65 -2747 -60
rect -2703 -70 -2699 -26
rect -2795 -74 -2699 -70
rect -2795 -85 -2791 -74
rect -2731 -85 -2727 -74
rect -2823 -89 -2818 -85
rect -2759 -89 -2754 -85
rect -2917 -106 -2913 -89
rect -2883 -106 -2879 -89
rect -2850 -106 -2846 -89
rect -2786 -106 -2782 -89
rect -2924 -121 -2767 -106
rect -2998 -209 -2772 -198
rect -2998 -424 -2991 -209
rect -2936 -210 -2772 -209
rect -2918 -243 -2914 -210
rect -2884 -243 -2880 -210
rect -2851 -243 -2847 -210
rect -2819 -243 -2815 -210
rect -2764 -224 -2699 -218
rect -2764 -243 -2760 -224
rect -2732 -243 -2728 -224
rect -2923 -287 -2915 -281
rect -2895 -332 -2891 -247
rect -2861 -282 -2857 -247
rect -2828 -271 -2824 -247
rect -2796 -271 -2792 -247
rect -2787 -271 -2783 -247
rect -2755 -271 -2751 -247
rect -2828 -275 -2751 -271
rect -2886 -288 -2879 -282
rect -2861 -288 -2812 -282
rect -2861 -332 -2857 -288
rect -2704 -295 -2699 -224
rect -2660 -295 -2649 -150
rect -2612 -295 -2605 -294
rect -2705 -300 -2605 -295
rect -2752 -312 -2748 -307
rect -2704 -317 -2699 -300
rect -2660 -301 -2649 -300
rect -2796 -321 -2699 -317
rect -2612 -320 -2605 -300
rect -2796 -332 -2792 -321
rect -2732 -332 -2728 -321
rect -2824 -336 -2819 -332
rect -2760 -336 -2755 -332
rect -2918 -353 -2914 -336
rect -2884 -353 -2880 -336
rect -2851 -353 -2847 -336
rect -2787 -352 -2783 -336
rect -2590 -347 -2587 -26
rect -2521 -262 -2512 36
rect -2169 -1 -2157 74
rect -2487 -146 -2210 -137
rect -2571 -271 -2269 -262
rect -2571 -277 -2295 -271
rect -2564 -289 -2560 -277
rect -2520 -289 -2516 -277
rect -2476 -289 -2472 -277
rect -2432 -289 -2428 -277
rect -2388 -289 -2384 -277
rect -2344 -289 -2340 -277
rect -2528 -304 -2524 -293
rect -2484 -304 -2480 -293
rect -2440 -304 -2436 -293
rect -2396 -304 -2392 -293
rect -2352 -304 -2348 -293
rect -2528 -308 -2348 -304
rect -2352 -342 -2343 -308
rect -2308 -339 -2304 -293
rect -2277 -317 -2270 -271
rect -2172 -330 -2157 -1
rect -2029 -286 -2007 -148
rect -2009 -304 -2007 -286
rect -1854 -330 -1839 60
rect -2566 -347 -2557 -346
rect -2788 -353 -2628 -352
rect -2918 -368 -2628 -353
rect -2590 -355 -2557 -347
rect -2516 -356 -2512 -347
rect -2467 -357 -2464 -348
rect -2426 -357 -2421 -348
rect -2382 -358 -2377 -350
rect -2386 -359 -2377 -358
rect -2352 -351 -2336 -342
rect -2308 -351 -2296 -339
rect -2172 -342 -1835 -330
rect -2788 -369 -2628 -368
rect -2636 -411 -2628 -369
rect -2352 -392 -2348 -351
rect -2308 -392 -2304 -351
rect -2524 -396 -2520 -392
rect -2480 -396 -2476 -392
rect -2436 -396 -2432 -392
rect -2392 -396 -2388 -392
rect -2564 -410 -2560 -396
rect -2344 -410 -2340 -396
rect -2567 -411 -2291 -410
rect -2998 -435 -2768 -424
rect -2636 -425 -2291 -411
rect -2998 -478 -2991 -435
rect -2932 -436 -2768 -435
rect -2914 -469 -2910 -436
rect -2880 -469 -2876 -436
rect -2847 -469 -2843 -436
rect -2815 -469 -2811 -436
rect -2760 -450 -2695 -444
rect -2760 -469 -2756 -450
rect -2728 -469 -2724 -450
rect -2999 -631 -2991 -478
rect -2919 -513 -2911 -507
rect -2891 -558 -2887 -473
rect -2857 -508 -2853 -473
rect -2824 -497 -2820 -473
rect -2792 -497 -2788 -473
rect -2700 -453 -2695 -450
rect -2700 -459 -2476 -453
rect -2783 -497 -2779 -473
rect -2751 -497 -2747 -473
rect -2824 -501 -2747 -497
rect -2882 -514 -2875 -508
rect -2857 -514 -2808 -508
rect -2857 -558 -2853 -514
rect -2748 -538 -2744 -533
rect -2700 -543 -2695 -459
rect -2792 -547 -2695 -543
rect -2792 -558 -2788 -547
rect -2728 -558 -2724 -547
rect -2820 -562 -2815 -558
rect -2756 -562 -2751 -558
rect -2914 -579 -2910 -562
rect -2880 -579 -2876 -562
rect -2847 -579 -2843 -562
rect -2783 -579 -2779 -562
rect -2912 -594 -2764 -579
rect -2435 -627 -2423 -460
rect -2172 -613 -2157 -342
rect -1854 -343 -1839 -342
rect -2172 -627 -2158 -613
rect -2999 -642 -2771 -631
rect -2988 -868 -2977 -642
rect -2935 -643 -2771 -642
rect -2917 -676 -2913 -643
rect -2883 -676 -2879 -643
rect -2850 -676 -2846 -643
rect -2818 -676 -2814 -643
rect -2435 -644 -2158 -627
rect -2763 -657 -2697 -651
rect -2763 -676 -2759 -657
rect -2731 -676 -2727 -657
rect -2922 -720 -2914 -714
rect -2894 -765 -2890 -680
rect -2860 -715 -2856 -680
rect -2827 -704 -2823 -680
rect -2795 -704 -2791 -680
rect -2786 -704 -2782 -680
rect -2754 -704 -2750 -680
rect -2827 -708 -2750 -704
rect -2703 -696 -2698 -657
rect -2435 -696 -2423 -644
rect -2172 -645 -2158 -644
rect -2703 -697 -2423 -696
rect -2703 -705 -2674 -697
rect -2666 -705 -2423 -697
rect -2885 -721 -2878 -715
rect -2860 -721 -2811 -715
rect -2860 -765 -2856 -721
rect -2751 -745 -2747 -740
rect -2703 -750 -2698 -705
rect -2795 -754 -2697 -750
rect -2795 -765 -2791 -754
rect -2731 -765 -2727 -754
rect -2823 -769 -2818 -765
rect -2759 -769 -2754 -765
rect -2917 -785 -2913 -769
rect -2914 -786 -2913 -785
rect -2883 -786 -2879 -769
rect -2850 -786 -2846 -769
rect -2786 -786 -2782 -769
rect -2914 -792 -2767 -786
rect -1441 -792 -1436 279
rect -2914 -799 -1436 -792
rect -2260 -831 -1471 -819
rect -2464 -857 -2458 -854
rect -2334 -857 -2328 -856
rect -2465 -862 -2328 -857
rect -2464 -868 -2458 -862
rect -2334 -867 -2328 -862
rect -2083 -858 -2076 -857
rect -1957 -858 -1950 -857
rect -2083 -861 -1949 -858
rect -2083 -867 -2076 -861
rect -1957 -867 -1950 -861
rect -2988 -869 -2891 -868
rect -2988 -870 -2794 -869
rect -2711 -870 -2439 -868
rect -2988 -876 -2439 -870
rect -2942 -993 -2934 -876
rect -2890 -885 -2885 -876
rect -2859 -885 -2854 -876
rect -2826 -885 -2821 -876
rect -2711 -877 -2439 -876
rect -2339 -874 -2067 -867
rect -1965 -874 -1689 -867
rect -2711 -883 -2435 -877
rect -2339 -882 -2063 -874
rect -1965 -877 -1565 -874
rect -1965 -882 -1689 -877
rect -2871 -914 -2866 -890
rect -2840 -914 -2835 -890
rect -2871 -920 -2821 -914
rect -2807 -917 -2802 -890
rect -2704 -895 -2700 -883
rect -2660 -895 -2656 -883
rect -2616 -895 -2612 -883
rect -2572 -895 -2568 -883
rect -2528 -895 -2524 -883
rect -2484 -895 -2480 -883
rect -2332 -894 -2328 -882
rect -2288 -894 -2284 -882
rect -2244 -894 -2240 -882
rect -2200 -894 -2196 -882
rect -2156 -894 -2152 -882
rect -2112 -894 -2108 -882
rect -1958 -894 -1954 -882
rect -1914 -894 -1910 -882
rect -1870 -894 -1866 -882
rect -1826 -894 -1822 -882
rect -1782 -894 -1778 -882
rect -1738 -894 -1734 -882
rect -2668 -910 -2664 -899
rect -2624 -910 -2620 -899
rect -2580 -910 -2576 -899
rect -2536 -910 -2532 -899
rect -2492 -910 -2488 -899
rect -2668 -914 -2488 -910
rect -2807 -918 -2759 -917
rect -2921 -933 -2884 -928
rect -2859 -933 -2853 -928
rect -2921 -975 -2916 -933
rect -2840 -943 -2835 -920
rect -2807 -922 -2758 -918
rect -2807 -943 -2802 -922
rect -2866 -948 -2859 -943
rect -2890 -952 -2885 -948
rect -2826 -952 -2821 -948
rect -2889 -959 -2789 -952
rect -2921 -978 -2769 -975
rect -2888 -993 -2798 -989
rect -2942 -999 -2798 -993
rect -2870 -1011 -2866 -999
rect -2857 -1036 -2852 -1032
rect -2822 -1033 -2818 -1015
rect -2774 -1033 -2769 -978
rect -2822 -1039 -2769 -1033
rect -2822 -1049 -2818 -1039
rect -2870 -1078 -2866 -1053
rect -2881 -1088 -2804 -1078
rect -2762 -1220 -2758 -922
rect -2492 -948 -2483 -914
rect -2730 -961 -2697 -952
rect -2661 -954 -2652 -953
rect -2730 -1148 -2726 -961
rect -2657 -962 -2652 -954
rect -2613 -963 -2604 -954
rect -2564 -963 -2561 -954
rect -2522 -965 -2517 -956
rect -2492 -957 -2476 -948
rect -2448 -956 -2444 -899
rect -2296 -909 -2292 -898
rect -2252 -909 -2248 -898
rect -2208 -909 -2204 -898
rect -2164 -909 -2160 -898
rect -2120 -909 -2116 -898
rect -2296 -913 -2116 -909
rect -2120 -947 -2111 -913
rect -2076 -943 -2072 -898
rect -1922 -909 -1918 -898
rect -1878 -909 -1874 -898
rect -1834 -909 -1830 -898
rect -1790 -909 -1786 -898
rect -1746 -909 -1742 -898
rect -1922 -913 -1742 -909
rect -2448 -957 -2436 -956
rect -2492 -998 -2488 -957
rect -2448 -998 -2444 -957
rect -2664 -1002 -2660 -998
rect -2620 -1002 -2616 -998
rect -2576 -1002 -2572 -998
rect -2532 -1002 -2528 -998
rect -2367 -961 -2325 -951
rect -2285 -961 -2280 -952
rect -2704 -1012 -2700 -1002
rect -2706 -1017 -2700 -1012
rect -2484 -1016 -2480 -1002
rect -2697 -1017 -2431 -1016
rect -2706 -1022 -2443 -1017
rect -2714 -1024 -2443 -1022
rect -2715 -1030 -2443 -1024
rect -2715 -1073 -2707 -1030
rect -2697 -1031 -2443 -1030
rect -2687 -1044 -2397 -1035
rect -2367 -1042 -2362 -961
rect -2235 -962 -2232 -953
rect -2198 -962 -2189 -953
rect -2147 -964 -2145 -955
rect -2120 -956 -2104 -947
rect -2120 -997 -2116 -956
rect -2076 -957 -2025 -943
rect -1746 -947 -1737 -913
rect -1702 -944 -1698 -898
rect -1573 -924 -1566 -877
rect -1510 -924 -1324 -923
rect -1573 -927 -1324 -924
rect -1510 -931 -1324 -927
rect -1702 -947 -1690 -944
rect -1498 -946 -1494 -931
rect -1365 -946 -1361 -931
rect -2076 -997 -2072 -957
rect -2292 -1001 -2288 -997
rect -2248 -1001 -2244 -997
rect -2204 -1001 -2200 -997
rect -2160 -1001 -2156 -997
rect -2332 -1013 -2328 -1001
rect -2112 -1015 -2108 -1001
rect -2327 -1028 -2066 -1015
rect -2335 -1030 -2059 -1028
rect -2171 -1042 -2168 -1041
rect -2687 -1045 -2593 -1044
rect -2673 -1057 -2669 -1045
rect -2625 -1078 -2621 -1061
rect -2405 -1059 -2398 -1044
rect -2367 -1048 -2168 -1042
rect -2405 -1069 -2199 -1059
rect -2186 -1069 -2185 -1059
rect -2405 -1070 -2398 -1069
rect -2660 -1082 -2655 -1078
rect -2715 -1126 -2704 -1090
rect -2625 -1085 -2570 -1078
rect -2265 -1081 -2261 -1069
rect -2625 -1095 -2621 -1085
rect -2673 -1124 -2669 -1099
rect -2680 -1126 -2608 -1124
rect -2715 -1133 -2608 -1126
rect -2680 -1134 -2594 -1133
rect -2577 -1148 -2570 -1085
rect -2252 -1106 -2247 -1102
rect -2217 -1103 -2213 -1085
rect -2171 -1103 -2168 -1048
rect -2217 -1109 -2166 -1103
rect -2217 -1119 -2213 -1109
rect -2265 -1148 -2261 -1123
rect -2730 -1151 -2570 -1148
rect -2577 -1152 -2570 -1151
rect -2275 -1158 -2199 -1148
rect -2035 -1184 -2025 -957
rect -1988 -960 -1951 -955
rect -1988 -1046 -1981 -960
rect -1911 -961 -1906 -952
rect -1861 -962 -1858 -953
rect -1819 -962 -1815 -953
rect -1789 -955 -1773 -953
rect -1789 -964 -1771 -955
rect -1746 -956 -1730 -947
rect -1702 -956 -1552 -947
rect -1469 -950 -1464 -946
rect -1435 -950 -1431 -946
rect -1402 -950 -1398 -946
rect -1746 -997 -1742 -956
rect -1702 -997 -1698 -956
rect -1564 -976 -1554 -956
rect -1564 -979 -1392 -976
rect -1494 -991 -1490 -990
rect -1918 -1001 -1914 -997
rect -1874 -1001 -1870 -997
rect -1830 -1001 -1826 -997
rect -1786 -1001 -1782 -997
rect -1529 -994 -1490 -991
rect -1529 -996 -1491 -994
rect -1458 -995 -1455 -991
rect -1395 -990 -1392 -979
rect -1423 -996 -1422 -992
rect -1958 -1015 -1954 -1001
rect -1738 -1015 -1734 -1001
rect -1961 -1016 -1697 -1015
rect -1951 -1029 -1697 -1016
rect -1951 -1030 -1685 -1029
rect -1988 -1050 -1732 -1046
rect -1988 -1052 -1733 -1050
rect -1848 -1068 -1758 -1058
rect -1838 -1080 -1834 -1068
rect -1825 -1105 -1820 -1101
rect -1790 -1102 -1786 -1084
rect -1790 -1104 -1782 -1102
rect -1736 -1104 -1733 -1052
rect -1790 -1108 -1733 -1104
rect -1790 -1118 -1786 -1108
rect -1736 -1109 -1733 -1108
rect -1838 -1147 -1834 -1122
rect -1848 -1157 -1771 -1147
rect -2035 -1199 -1594 -1184
rect -1529 -1220 -1523 -996
rect -1373 -991 -1369 -950
rect -1340 -991 -1336 -950
rect -1390 -997 -1389 -993
rect -1373 -995 -1357 -991
rect -1340 -995 -1327 -991
rect -1373 -1007 -1369 -995
rect -1473 -1011 -1369 -1007
rect -1473 -1028 -1469 -1011
rect -1439 -1028 -1435 -1011
rect -1406 -1028 -1402 -1011
rect -1373 -1028 -1369 -1011
rect -1340 -1028 -1336 -995
rect -1498 -1037 -1494 -1032
rect -1464 -1040 -1460 -1032
rect -1431 -1040 -1427 -1032
rect -1398 -1040 -1394 -1032
rect -1365 -1040 -1361 -1032
rect -1492 -1048 -1315 -1040
rect -2762 -1226 -1521 -1220
<< m2contact >>
rect -2829 541 -2819 549
rect -2647 537 -2637 545
rect -2276 501 -2270 507
rect -2576 495 -2567 501
rect -2053 500 -2043 507
rect -2838 456 -2826 463
rect -2091 344 -2084 353
rect -1512 332 -1507 339
rect -2480 290 -2470 299
rect -2773 263 -2760 274
rect -2724 264 -2712 273
rect -2628 263 -2618 272
rect -2581 261 -2571 270
rect -2495 269 -2488 280
rect -2376 266 -2370 272
rect -2332 265 -2325 271
rect -2289 261 -2279 273
rect -2200 262 -2191 269
rect -2110 269 -2101 280
rect -1999 265 -1987 274
rect -1954 264 -1943 273
rect -1905 263 -1894 274
rect -1859 263 -1851 272
rect -1729 270 -1718 280
rect -2943 185 -2931 192
rect -2837 186 -2825 193
rect -2797 201 -2792 216
rect -1482 329 -1476 339
rect -1447 330 -1441 336
rect -1455 267 -1445 274
rect -2777 72 -2764 83
rect -2991 37 -2982 48
rect -2890 -65 -2882 -60
rect -2758 -65 -2751 -60
rect -2945 -122 -2924 -105
rect -2661 -150 -2644 -131
rect -2891 -312 -2883 -307
rect -2759 -312 -2752 -307
rect -2612 -336 -2605 -320
rect -2937 -368 -2918 -352
rect -2500 -146 -2487 -135
rect -2210 -148 -2193 -131
rect -2277 -331 -2269 -317
rect -1854 60 -1839 80
rect -2030 -148 -2007 -134
rect -2029 -304 -2009 -286
rect -2528 -356 -2516 -346
rect -2476 -358 -2467 -347
rect -2435 -358 -2426 -348
rect -2390 -358 -2382 -344
rect -2476 -459 -2466 -445
rect -2887 -538 -2879 -533
rect -2755 -538 -2748 -533
rect -2436 -460 -2422 -442
rect -2931 -595 -2912 -579
rect -2674 -705 -2666 -697
rect -2890 -745 -2882 -740
rect -2758 -745 -2751 -740
rect -2933 -799 -2914 -785
rect -2277 -831 -2260 -812
rect -1471 -831 -1460 -819
rect -2439 -877 -2431 -868
rect -2067 -874 -2055 -867
rect -2896 -959 -2889 -952
rect -2798 -1000 -2787 -989
rect -2890 -1090 -2881 -1078
rect -2804 -1092 -2790 -1077
rect -2665 -962 -2657 -954
rect -2572 -963 -2564 -954
rect -2530 -965 -2522 -956
rect -2444 -956 -2430 -945
rect -2294 -961 -2285 -952
rect -2443 -1032 -2429 -1017
rect -2698 -1046 -2687 -1035
rect -2248 -962 -2235 -953
rect -2157 -964 -2147 -955
rect -2341 -1028 -2327 -1013
rect -2066 -1028 -2052 -1013
rect -2720 -1090 -2704 -1073
rect -2199 -1069 -2186 -1059
rect -2608 -1133 -2594 -1118
rect -2289 -1163 -2275 -1148
rect -2199 -1159 -2185 -1144
rect -1924 -961 -1911 -952
rect -1874 -962 -1861 -953
rect -1832 -962 -1819 -953
rect -1463 -995 -1458 -988
rect -1428 -996 -1423 -989
rect -1965 -1031 -1951 -1016
rect -1697 -1029 -1683 -1014
rect -1861 -1068 -1848 -1058
rect -1862 -1158 -1848 -1143
rect -1771 -1160 -1757 -1145
rect -1594 -1207 -1564 -1174
rect -1395 -997 -1390 -990
rect -1506 -1052 -1492 -1037
<< metal2 >>
rect -2989 604 -2720 606
rect -2991 593 -2720 604
rect -2991 48 -2984 593
rect -2725 589 -2720 593
rect -2726 581 -2720 589
rect -2726 545 -2721 581
rect -2819 541 -2647 545
rect -2567 495 -2520 500
rect -2575 494 -2520 495
rect -2833 208 -2829 456
rect -2525 409 -2520 494
rect -2273 442 -2270 501
rect -2043 501 -2011 506
rect -2402 437 -2270 442
rect -2724 403 -2520 409
rect -2438 408 -2431 410
rect -2774 263 -2773 268
rect -2724 273 -2719 403
rect -2579 298 -2575 299
rect -2624 294 -2480 298
rect -2624 272 -2620 294
rect -2579 270 -2575 294
rect -2774 242 -2767 263
rect -2438 274 -2431 395
rect -2488 269 -2431 274
rect -2495 268 -2431 269
rect -2402 270 -2399 437
rect -2089 294 -2084 344
rect -2200 287 -2084 294
rect -2402 266 -2376 270
rect -2332 242 -2329 265
rect -2774 239 -2329 242
rect -2200 269 -2196 287
rect -2015 272 -2011 501
rect -1631 350 -1623 395
rect -1631 342 -1508 350
rect -1512 339 -1508 342
rect -2101 269 -2063 272
rect -2200 261 -2196 262
rect -2833 205 -2797 208
rect -2957 192 -2938 195
rect -2833 193 -2829 205
rect -2957 185 -2943 192
rect -2957 184 -2938 185
rect -2957 -105 -2951 184
rect -2774 83 -2767 239
rect -2289 162 -2281 261
rect -2294 161 -2281 162
rect -2475 157 -2281 161
rect -2068 159 -2064 269
rect -2015 268 -1999 272
rect -2475 21 -2469 157
rect -2068 156 -1986 159
rect -2882 -65 -2758 -60
rect -2957 -119 -2945 -105
rect -2955 -122 -2945 -119
rect -2955 -132 -2934 -122
rect -2954 -358 -2947 -132
rect -2644 -146 -2500 -139
rect -2644 -147 -2487 -146
rect -2475 -222 -2468 21
rect -2193 -148 -2030 -138
rect -1954 -138 -1945 264
rect -1718 270 -1636 274
rect -1481 271 -1477 329
rect -1447 274 -1444 330
rect -1720 269 -1636 270
rect -2007 -148 -1944 -138
rect -1903 -222 -1896 263
rect -1854 80 -1851 263
rect -1643 234 -1637 269
rect -1500 268 -1477 271
rect -1643 228 -1545 234
rect -1500 163 -1494 268
rect -1445 271 -1444 274
rect -1455 235 -1449 267
rect -2475 -231 -1889 -222
rect -2883 -312 -2759 -307
rect -2605 -336 -2521 -331
rect -2612 -337 -2521 -336
rect -2528 -346 -2521 -337
rect -2954 -367 -2937 -358
rect -2954 -581 -2947 -367
rect -2475 -347 -2468 -231
rect -1903 -233 -1896 -231
rect -2390 -331 -2277 -324
rect -2390 -335 -2269 -331
rect -2390 -344 -2382 -335
rect -2476 -445 -2469 -358
rect -2432 -442 -2428 -358
rect -2477 -459 -2476 -446
rect -2879 -538 -2755 -533
rect -2954 -586 -2942 -581
rect -2954 -595 -2931 -586
rect -2954 -793 -2947 -595
rect -2882 -745 -2758 -740
rect -2954 -799 -2933 -793
rect -2954 -808 -2943 -799
rect -2954 -1084 -2947 -808
rect -2670 -951 -2667 -705
rect -2477 -759 -2471 -459
rect -2025 -736 -2009 -304
rect -2025 -743 -2008 -736
rect -2025 -750 -1826 -743
rect -2023 -752 -1826 -750
rect -2477 -761 -2270 -759
rect -2248 -761 -2243 -760
rect -2477 -764 -2241 -761
rect -2476 -766 -2241 -764
rect -2275 -767 -2241 -766
rect -2403 -822 -2396 -820
rect -2403 -828 -2277 -822
rect -2431 -877 -2424 -871
rect -2428 -932 -2424 -877
rect -2572 -935 -2424 -932
rect -2910 -959 -2896 -954
rect -2670 -954 -2664 -951
rect -2572 -954 -2566 -935
rect -2910 -960 -2893 -959
rect -2910 -1084 -2901 -960
rect -2670 -962 -2665 -954
rect -2669 -980 -2663 -962
rect -2529 -956 -2523 -935
rect -2428 -936 -2424 -935
rect -2403 -950 -2396 -828
rect -2248 -845 -2243 -767
rect -2248 -851 -1861 -845
rect -2430 -956 -2395 -950
rect -2248 -953 -2243 -851
rect -2059 -932 -2056 -874
rect -2157 -936 -2056 -932
rect -2292 -980 -2289 -961
rect -2157 -955 -2154 -936
rect -1925 -961 -1924 -957
rect -1873 -953 -1865 -851
rect -1832 -953 -1826 -752
rect -1925 -980 -1918 -961
rect -1832 -963 -1826 -962
rect -2669 -984 -1917 -980
rect -1463 -988 -1460 -831
rect -2745 -991 -2742 -990
rect -2787 -998 -2742 -991
rect -2745 -1037 -2742 -998
rect -1430 -996 -1428 -989
rect -2429 -1028 -2341 -1018
rect -2052 -1023 -1965 -1020
rect -1683 -1028 -1512 -1022
rect -2745 -1044 -2698 -1037
rect -1519 -1041 -1513 -1028
rect -1519 -1049 -1506 -1041
rect -2186 -1068 -1861 -1061
rect -2954 -1089 -2890 -1084
rect -2954 -1093 -2947 -1089
rect -2790 -1088 -2720 -1079
rect -2594 -1131 -2307 -1127
rect -2320 -1150 -2314 -1131
rect -2320 -1158 -2289 -1150
rect -2185 -1158 -1862 -1151
rect -2185 -1159 -1856 -1158
rect -1519 -1147 -1513 -1049
rect -1757 -1154 -1511 -1147
rect -1430 -1186 -1424 -996
rect -1564 -1197 -1415 -1186
<< m3contact >>
rect -2438 395 -2428 408
rect -1633 395 -1622 404
rect -1986 156 -1978 163
rect -1545 228 -1534 238
rect -1455 228 -1445 235
rect -1500 156 -1494 163
<< metal3 >>
rect -2428 395 -1633 404
rect -1534 228 -1455 234
rect -1978 156 -1500 161
<< labels >>
rlabel metal1 -2305 -345 -2305 -345 1 node_c2
rlabel metal1 -2845 -118 -2845 -118 1 gnd
rlabel metal1 -2930 41 -2930 41 1 vdd
rlabel metal1 -2882 -718 -2882 -718 1 node_b3
rlabel metal1 -2920 -717 -2920 -717 1 node_a3
rlabel metal1 -2878 -512 -2878 -512 1 node_b2
rlabel metal1 -2915 -511 -2915 -511 1 node_a2
rlabel metal1 -2884 -285 -2884 -285 1 node_b1
rlabel metal1 -2920 -284 -2920 -284 1 node_a1
rlabel metal1 -2882 -37 -2882 -37 1 node_b0
rlabel metal1 -2920 -39 -2920 -39 1 node_a0
rlabel metal1 -2714 225 -2714 225 1 node_x
rlabel metal1 -2332 225 -2332 225 1 node_x
rlabel metal1 -1950 225 -1950 225 1 node_x
rlabel metal1 -2882 504 -2882 504 1 node_b3
rlabel metal1 -2612 500 -2612 500 1 node_b2
rlabel metal1 -2357 506 -2357 506 1 node_b1
rlabel metal1 -2090 505 -2090 505 1 node_b0
rlabel metal1 -2901 215 -2901 215 1 node_a3
rlabel metal1 -2661 269 -2661 269 1 node_a2
rlabel metal1 -2235 267 -2235 267 1 node_a1
rlabel metal1 -1809 262 -1809 262 1 node_a0
rlabel metal1 -1383 334 -1383 334 1 node_c1
rlabel metal1 -2856 -1034 -2856 -1034 1 node_a3
rlabel metal1 -2857 -930 -2857 -930 1 node_b3
rlabel metal1 -2659 -1081 -2659 -1081 1 node_a2
rlabel metal1 -2610 -960 -2610 -960 1 node_b2
rlabel metal1 -2249 -1104 -2249 -1104 1 node_a1
rlabel metal1 -2194 -959 -2194 -959 1 node_b1
rlabel metal1 -1824 -1104 -1824 -1104 1 node_a0
rlabel metal1 -1782 -958 -1782 -958 1 node_b0
rlabel metal1 -1332 -993 -1332 -993 1 node_c3
<< end >>
