magic
tech scmos
timestamp 1699186971
<< nwell >>
rect -565 470 -377 509
<< ntransistor >>
rect -550 412 -547 419
rect -521 412 -519 419
rect -490 412 -487 419
rect -461 412 -458 419
rect -432 412 -429 419
rect -402 412 -399 419
<< ptransistor >>
rect -550 484 -547 491
rect -521 484 -519 491
rect -490 484 -487 491
rect -461 484 -458 491
rect -432 484 -429 491
rect -402 484 -399 491
<< ndiffusion >>
rect -555 415 -550 419
rect -559 412 -550 415
rect -547 415 -538 419
rect -547 412 -534 415
rect -526 415 -521 419
rect -530 412 -521 415
rect -519 415 -509 419
rect -519 412 -505 415
rect -497 415 -490 419
rect -501 412 -490 415
rect -487 415 -480 419
rect -487 412 -476 415
rect -468 415 -461 419
rect -472 412 -461 415
rect -458 415 -451 419
rect -458 412 -447 415
rect -439 415 -432 419
rect -443 412 -432 415
rect -429 415 -422 419
rect -429 412 -418 415
rect -410 415 -402 419
rect -414 412 -402 415
rect -399 415 -393 419
rect -399 412 -389 415
<< pdiffusion >>
rect -555 487 -550 491
rect -559 484 -550 487
rect -547 487 -538 491
rect -547 484 -534 487
rect -526 487 -521 491
rect -530 484 -521 487
rect -519 487 -509 491
rect -519 484 -505 487
rect -497 487 -490 491
rect -501 484 -490 487
rect -487 487 -480 491
rect -487 484 -476 487
rect -468 487 -461 491
rect -472 484 -461 487
rect -458 487 -451 491
rect -458 484 -447 487
rect -439 487 -432 491
rect -443 484 -432 487
rect -429 487 -422 491
rect -429 484 -418 487
rect -410 487 -402 491
rect -414 484 -402 487
rect -399 487 -393 491
rect -399 484 -389 487
<< ndcontact >>
rect -559 415 -555 419
rect -538 415 -534 419
rect -530 415 -526 419
rect -509 415 -505 419
rect -501 415 -497 419
rect -480 415 -476 419
rect -472 415 -468 419
rect -451 415 -447 419
rect -443 415 -439 419
rect -422 415 -418 419
rect -414 415 -410 419
rect -393 415 -389 419
<< pdcontact >>
rect -559 487 -555 491
rect -538 487 -534 491
rect -530 487 -526 491
rect -509 487 -505 491
rect -501 487 -497 491
rect -480 487 -476 491
rect -472 487 -468 491
rect -451 487 -447 491
rect -443 487 -439 491
rect -422 487 -418 491
rect -414 487 -410 491
rect -393 487 -389 491
<< polysilicon >>
rect -550 497 -487 499
rect -550 491 -547 497
rect -521 491 -519 494
rect -490 491 -487 497
rect -461 491 -458 495
rect -432 491 -429 495
rect -402 491 -399 495
rect -550 419 -547 484
rect -521 419 -519 484
rect -490 419 -487 484
rect -461 419 -458 484
rect -439 457 -436 462
rect -432 419 -429 484
rect -402 419 -399 484
rect -550 407 -547 412
rect -521 400 -519 412
rect -490 409 -487 412
rect -461 400 -458 412
rect -432 407 -429 412
rect -402 407 -399 412
rect -521 397 -458 400
<< polycontact >>
rect -555 448 -550 453
rect -526 447 -521 452
rect -436 457 -432 462
rect -407 430 -402 436
<< metal1 >>
rect -565 510 -377 517
rect -559 491 -555 510
rect -530 491 -526 510
rect -501 491 -497 510
rect -472 491 -468 510
rect -451 496 -410 500
rect -451 491 -447 496
rect -443 491 -439 496
rect -414 491 -410 496
rect -558 448 -555 453
rect -538 419 -534 487
rect -529 447 -526 452
rect -509 436 -505 487
rect -480 480 -476 487
rect -451 480 -447 487
rect -480 477 -447 480
rect -422 480 -418 487
rect -393 480 -389 487
rect -422 477 -389 480
rect -444 458 -436 462
rect -439 457 -436 458
rect -393 454 -389 477
rect -393 444 -385 454
rect -509 431 -407 436
rect -509 419 -505 431
rect -411 430 -407 431
rect -393 427 -389 444
rect -451 419 -447 420
rect -393 419 -389 422
rect -476 415 -472 419
rect -418 415 -414 419
rect -559 411 -555 415
rect -530 411 -526 415
rect -501 411 -497 415
rect -443 411 -439 415
rect -562 404 -374 411
<< m2contact >>
rect -534 458 -528 463
rect -449 458 -444 463
rect -451 420 -446 425
rect -394 422 -389 427
<< metal2 >>
rect -528 458 -449 462
rect -446 422 -394 425
<< labels >>
rlabel metal1 -519 513 -519 513 5 vdd
rlabel metal1 -557 450 -557 450 1 node_a
rlabel metal1 -528 448 -528 448 1 node_b
rlabel metal1 -537 460 -537 460 1 node_anot
rlabel metal1 -506 435 -506 435 1 node_bnot
rlabel metal1 -500 409 -500 409 1 gnd
rlabel metal1 -389 449 -389 449 1 node_out
rlabel metal1 -432 497 -432 497 1 node_x
rlabel metal1 -474 417 -474 417 1 node_y
rlabel metal1 -417 417 -417 417 1 node_z
<< end >>
