magic
tech scmos
timestamp 1700159819
<< nwell >>
rect -840 246 -652 285
rect -622 246 -434 285
rect -389 248 -201 287
rect -129 249 59 288
rect -811 48 -623 87
rect -584 48 -484 78
rect -411 34 -341 50
rect -185 45 3 84
rect 42 45 142 75
rect 215 31 285 47
rect 415 45 603 84
rect 642 45 742 75
rect 1018 48 1206 87
rect 1245 48 1345 78
rect 815 31 885 47
rect 1418 34 1488 50
rect -568 -91 -468 -61
rect 58 -94 158 -64
rect 658 -94 758 -64
rect 1261 -91 1361 -61
rect -801 -208 -613 -169
rect -175 -211 13 -172
rect 425 -211 613 -172
rect 1028 -208 1216 -169
<< ntransistor >>
rect -825 188 -822 195
rect -796 188 -794 195
rect -765 188 -762 195
rect -736 188 -733 195
rect -707 188 -704 195
rect -677 188 -674 195
rect -607 188 -604 195
rect -578 188 -576 195
rect -547 188 -544 195
rect -518 188 -515 195
rect -489 188 -486 195
rect -459 188 -456 195
rect -374 190 -371 197
rect -345 190 -343 197
rect -314 190 -311 197
rect -285 190 -282 197
rect -256 190 -253 197
rect -226 190 -223 197
rect -114 191 -111 198
rect -85 191 -83 198
rect -54 191 -51 198
rect -25 191 -22 198
rect 4 191 7 198
rect 34 191 37 198
rect -569 2 -565 11
rect -537 2 -533 11
rect -503 2 -499 11
rect -396 -1 -394 3
rect -378 -1 -376 3
rect -359 -1 -357 3
rect -796 -10 -793 -3
rect -767 -10 -765 -3
rect -736 -10 -733 -3
rect -707 -10 -704 -3
rect -678 -10 -675 -3
rect -648 -10 -645 -3
rect 57 -1 61 8
rect 89 -1 93 8
rect 123 -1 127 8
rect 230 -4 232 0
rect 248 -4 250 0
rect 267 -4 269 0
rect -170 -13 -167 -6
rect -141 -13 -139 -6
rect -110 -13 -107 -6
rect -81 -13 -78 -6
rect -52 -13 -49 -6
rect -22 -13 -19 -6
rect 657 -1 661 8
rect 689 -1 693 8
rect 723 -1 727 8
rect 830 -4 832 0
rect 848 -4 850 0
rect 867 -4 869 0
rect 1260 2 1264 11
rect 1292 2 1296 11
rect 1326 2 1330 11
rect 1433 -1 1435 3
rect 1451 -1 1453 3
rect 1470 -1 1472 3
rect 430 -13 433 -6
rect 459 -13 461 -6
rect 490 -13 493 -6
rect 519 -13 522 -6
rect 548 -13 551 -6
rect 578 -13 581 -6
rect 1033 -10 1036 -3
rect 1062 -10 1064 -3
rect 1093 -10 1096 -3
rect 1122 -10 1125 -3
rect 1151 -10 1154 -3
rect 1181 -10 1184 -3
rect -553 -137 -549 -128
rect -521 -137 -517 -128
rect -487 -137 -483 -128
rect 73 -140 77 -131
rect 105 -140 109 -131
rect 139 -140 143 -131
rect 673 -140 677 -131
rect 705 -140 709 -131
rect 739 -140 743 -131
rect 1276 -137 1280 -128
rect 1308 -137 1312 -128
rect 1342 -137 1346 -128
rect -786 -266 -783 -259
rect -757 -266 -755 -259
rect -726 -266 -723 -259
rect -697 -266 -694 -259
rect -668 -266 -665 -259
rect -638 -266 -635 -259
rect -160 -269 -157 -262
rect -131 -269 -129 -262
rect -100 -269 -97 -262
rect -71 -269 -68 -262
rect -42 -269 -39 -262
rect -12 -269 -9 -262
rect 440 -269 443 -262
rect 469 -269 471 -262
rect 500 -269 503 -262
rect 529 -269 532 -262
rect 558 -269 561 -262
rect 588 -269 591 -262
rect 1043 -266 1046 -259
rect 1072 -266 1074 -259
rect 1103 -266 1106 -259
rect 1132 -266 1135 -259
rect 1161 -266 1164 -259
rect 1191 -266 1194 -259
<< ptransistor >>
rect -825 260 -822 267
rect -796 260 -794 267
rect -765 260 -762 267
rect -736 260 -733 267
rect -707 260 -704 267
rect -677 260 -674 267
rect -607 260 -604 267
rect -578 260 -576 267
rect -547 260 -544 267
rect -518 260 -515 267
rect -489 260 -486 267
rect -459 260 -456 267
rect -374 262 -371 269
rect -345 262 -343 269
rect -314 262 -311 269
rect -285 262 -282 269
rect -256 262 -253 269
rect -226 262 -223 269
rect -114 263 -111 270
rect -85 263 -83 270
rect -54 263 -51 270
rect -25 263 -22 270
rect 4 263 7 270
rect 34 263 37 270
rect -796 62 -793 69
rect -767 62 -765 69
rect -736 62 -733 69
rect -707 62 -704 69
rect -678 62 -675 69
rect -648 62 -645 69
rect -569 60 -565 69
rect -537 60 -533 69
rect -503 60 -499 69
rect -170 59 -167 66
rect -141 59 -139 66
rect -110 59 -107 66
rect -81 59 -78 66
rect -52 59 -49 66
rect -22 59 -19 66
rect -396 40 -394 44
rect -378 40 -376 44
rect -359 40 -357 44
rect 57 57 61 66
rect 89 57 93 66
rect 123 57 127 66
rect 430 59 433 66
rect 459 59 461 66
rect 490 59 493 66
rect 519 59 522 66
rect 548 59 551 66
rect 578 59 581 66
rect 230 37 232 41
rect 248 37 250 41
rect 267 37 269 41
rect 657 57 661 66
rect 689 57 693 66
rect 723 57 727 66
rect 1033 62 1036 69
rect 1062 62 1064 69
rect 1093 62 1096 69
rect 1122 62 1125 69
rect 1151 62 1154 69
rect 1181 62 1184 69
rect 830 37 832 41
rect 848 37 850 41
rect 867 37 869 41
rect 1260 60 1264 69
rect 1292 60 1296 69
rect 1326 60 1330 69
rect 1433 40 1435 44
rect 1451 40 1453 44
rect 1470 40 1472 44
rect -553 -79 -549 -70
rect -521 -79 -517 -70
rect -487 -79 -483 -70
rect 73 -82 77 -73
rect 105 -82 109 -73
rect 139 -82 143 -73
rect 673 -82 677 -73
rect 705 -82 709 -73
rect 739 -82 743 -73
rect 1276 -79 1280 -70
rect 1308 -79 1312 -70
rect 1342 -79 1346 -70
rect -786 -194 -783 -187
rect -757 -194 -755 -187
rect -726 -194 -723 -187
rect -697 -194 -694 -187
rect -668 -194 -665 -187
rect -638 -194 -635 -187
rect -160 -197 -157 -190
rect -131 -197 -129 -190
rect -100 -197 -97 -190
rect -71 -197 -68 -190
rect -42 -197 -39 -190
rect -12 -197 -9 -190
rect 440 -197 443 -190
rect 469 -197 471 -190
rect 500 -197 503 -190
rect 529 -197 532 -190
rect 558 -197 561 -190
rect 588 -197 591 -190
rect 1043 -194 1046 -187
rect 1072 -194 1074 -187
rect 1103 -194 1106 -187
rect 1132 -194 1135 -187
rect 1161 -194 1164 -187
rect 1191 -194 1194 -187
<< ndiffusion >>
rect -830 191 -825 195
rect -834 188 -825 191
rect -822 191 -813 195
rect -822 188 -809 191
rect -801 191 -796 195
rect -805 188 -796 191
rect -794 191 -784 195
rect -794 188 -780 191
rect -772 191 -765 195
rect -776 188 -765 191
rect -762 191 -755 195
rect -762 188 -751 191
rect -743 191 -736 195
rect -747 188 -736 191
rect -733 191 -726 195
rect -733 188 -722 191
rect -714 191 -707 195
rect -718 188 -707 191
rect -704 191 -697 195
rect -704 188 -693 191
rect -685 191 -677 195
rect -689 188 -677 191
rect -674 191 -668 195
rect -674 188 -664 191
rect -612 191 -607 195
rect -616 188 -607 191
rect -604 191 -595 195
rect -604 188 -591 191
rect -583 191 -578 195
rect -587 188 -578 191
rect -576 191 -566 195
rect -576 188 -562 191
rect -554 191 -547 195
rect -558 188 -547 191
rect -544 191 -537 195
rect -544 188 -533 191
rect -525 191 -518 195
rect -529 188 -518 191
rect -515 191 -508 195
rect -515 188 -504 191
rect -496 191 -489 195
rect -500 188 -489 191
rect -486 191 -479 195
rect -486 188 -475 191
rect -467 191 -459 195
rect -471 188 -459 191
rect -456 191 -450 195
rect -456 188 -446 191
rect -379 193 -374 197
rect -383 190 -374 193
rect -371 193 -362 197
rect -371 190 -358 193
rect -350 193 -345 197
rect -354 190 -345 193
rect -343 193 -333 197
rect -343 190 -329 193
rect -321 193 -314 197
rect -325 190 -314 193
rect -311 193 -304 197
rect -311 190 -300 193
rect -292 193 -285 197
rect -296 190 -285 193
rect -282 193 -275 197
rect -282 190 -271 193
rect -263 193 -256 197
rect -267 190 -256 193
rect -253 193 -246 197
rect -253 190 -242 193
rect -234 193 -226 197
rect -238 190 -226 193
rect -223 193 -217 197
rect -223 190 -213 193
rect -119 194 -114 198
rect -123 191 -114 194
rect -111 194 -102 198
rect -111 191 -98 194
rect -90 194 -85 198
rect -94 191 -85 194
rect -83 194 -73 198
rect -83 191 -69 194
rect -61 194 -54 198
rect -65 191 -54 194
rect -51 194 -44 198
rect -51 191 -40 194
rect -32 194 -25 198
rect -36 191 -25 194
rect -22 194 -15 198
rect -22 191 -11 194
rect -3 194 4 198
rect -7 191 4 194
rect 7 194 14 198
rect 7 191 18 194
rect 26 194 34 198
rect 22 191 34 194
rect 37 194 43 198
rect 37 191 47 194
rect -573 6 -569 11
rect -578 2 -569 6
rect -565 6 -559 11
rect -565 2 -554 6
rect -542 6 -537 11
rect -547 2 -537 6
rect -533 6 -528 11
rect -533 2 -523 6
rect -509 6 -503 11
rect -514 2 -503 6
rect -499 6 -495 11
rect -499 2 -490 6
rect -398 -1 -396 3
rect -394 -1 -392 3
rect -380 -1 -378 3
rect -376 -1 -374 3
rect -361 -1 -359 3
rect -357 -1 -355 3
rect -801 -7 -796 -3
rect -805 -10 -796 -7
rect -793 -7 -784 -3
rect -793 -10 -780 -7
rect -772 -7 -767 -3
rect -776 -10 -767 -7
rect -765 -7 -755 -3
rect -765 -10 -751 -7
rect -743 -7 -736 -3
rect -747 -10 -736 -7
rect -733 -7 -726 -3
rect -733 -10 -722 -7
rect -714 -7 -707 -3
rect -718 -10 -707 -7
rect -704 -7 -697 -3
rect -704 -10 -693 -7
rect -685 -7 -678 -3
rect -689 -10 -678 -7
rect -675 -7 -668 -3
rect -675 -10 -664 -7
rect -656 -7 -648 -3
rect -660 -10 -648 -7
rect -645 -7 -639 -3
rect 53 3 57 8
rect 48 -1 57 3
rect 61 3 67 8
rect 61 -1 72 3
rect 84 3 89 8
rect 79 -1 89 3
rect 93 3 98 8
rect 93 -1 103 3
rect 117 3 123 8
rect 112 -1 123 3
rect 127 3 131 8
rect 127 -1 136 3
rect 228 -4 230 0
rect 232 -4 234 0
rect 246 -4 248 0
rect 250 -4 252 0
rect 265 -4 267 0
rect 269 -4 271 0
rect -645 -10 -635 -7
rect -175 -10 -170 -6
rect -179 -13 -170 -10
rect -167 -10 -158 -6
rect -167 -13 -154 -10
rect -146 -10 -141 -6
rect -150 -13 -141 -10
rect -139 -10 -129 -6
rect -139 -13 -125 -10
rect -117 -10 -110 -6
rect -121 -13 -110 -10
rect -107 -10 -100 -6
rect -107 -13 -96 -10
rect -88 -10 -81 -6
rect -92 -13 -81 -10
rect -78 -10 -71 -6
rect -78 -13 -67 -10
rect -59 -10 -52 -6
rect -63 -13 -52 -10
rect -49 -10 -42 -6
rect -49 -13 -38 -10
rect -30 -10 -22 -6
rect -34 -13 -22 -10
rect -19 -10 -13 -6
rect 653 3 657 8
rect 648 -1 657 3
rect 661 3 667 8
rect 661 -1 672 3
rect 684 3 689 8
rect 679 -1 689 3
rect 693 3 698 8
rect 693 -1 703 3
rect 717 3 723 8
rect 712 -1 723 3
rect 727 3 731 8
rect 727 -1 736 3
rect 828 -4 830 0
rect 832 -4 834 0
rect 846 -4 848 0
rect 850 -4 852 0
rect 865 -4 867 0
rect 869 -4 871 0
rect 1256 6 1260 11
rect 1251 2 1260 6
rect 1264 6 1270 11
rect 1264 2 1275 6
rect 1287 6 1292 11
rect 1282 2 1292 6
rect 1296 6 1301 11
rect 1296 2 1306 6
rect 1320 6 1326 11
rect 1315 2 1326 6
rect 1330 6 1334 11
rect 1330 2 1339 6
rect 1431 -1 1433 3
rect 1435 -1 1437 3
rect 1449 -1 1451 3
rect 1453 -1 1455 3
rect 1468 -1 1470 3
rect 1472 -1 1474 3
rect -19 -13 -9 -10
rect 425 -10 430 -6
rect 421 -13 430 -10
rect 433 -10 442 -6
rect 433 -13 446 -10
rect 454 -10 459 -6
rect 450 -13 459 -10
rect 461 -10 471 -6
rect 461 -13 475 -10
rect 483 -10 490 -6
rect 479 -13 490 -10
rect 493 -10 500 -6
rect 493 -13 504 -10
rect 512 -10 519 -6
rect 508 -13 519 -10
rect 522 -10 529 -6
rect 522 -13 533 -10
rect 541 -10 548 -6
rect 537 -13 548 -10
rect 551 -10 558 -6
rect 551 -13 562 -10
rect 570 -10 578 -6
rect 566 -13 578 -10
rect 581 -10 587 -6
rect 1028 -7 1033 -3
rect 1024 -10 1033 -7
rect 1036 -7 1045 -3
rect 1036 -10 1049 -7
rect 1057 -7 1062 -3
rect 1053 -10 1062 -7
rect 1064 -7 1074 -3
rect 1064 -10 1078 -7
rect 1086 -7 1093 -3
rect 1082 -9 1093 -7
rect 1085 -10 1093 -9
rect 1096 -7 1103 -3
rect 1096 -10 1107 -7
rect 1115 -7 1122 -3
rect 1111 -10 1122 -7
rect 1125 -7 1132 -3
rect 1125 -10 1136 -7
rect 1144 -7 1151 -3
rect 1140 -10 1151 -7
rect 1154 -7 1161 -3
rect 1154 -10 1165 -7
rect 1173 -7 1181 -3
rect 1169 -10 1181 -7
rect 1184 -7 1190 -3
rect 1184 -10 1194 -7
rect 581 -13 591 -10
rect -557 -133 -553 -128
rect -562 -137 -553 -133
rect -549 -133 -543 -128
rect -549 -137 -538 -133
rect -526 -133 -521 -128
rect -531 -137 -521 -133
rect -517 -133 -512 -128
rect -517 -137 -507 -133
rect -493 -133 -487 -128
rect -498 -137 -487 -133
rect -483 -133 -479 -128
rect -483 -137 -474 -133
rect 69 -136 73 -131
rect 64 -140 73 -136
rect 77 -136 83 -131
rect 77 -140 88 -136
rect 100 -136 105 -131
rect 95 -140 105 -136
rect 109 -136 114 -131
rect 109 -140 119 -136
rect 133 -136 139 -131
rect 128 -140 139 -136
rect 143 -136 147 -131
rect 143 -140 152 -136
rect 669 -136 673 -131
rect 664 -140 673 -136
rect 677 -136 683 -131
rect 677 -140 688 -136
rect 700 -136 705 -131
rect 695 -140 705 -136
rect 709 -136 714 -131
rect 709 -140 719 -136
rect 733 -136 739 -131
rect 728 -140 739 -136
rect 743 -136 747 -131
rect 743 -140 752 -136
rect 1272 -133 1276 -128
rect 1267 -137 1276 -133
rect 1280 -133 1286 -128
rect 1280 -137 1291 -133
rect 1303 -133 1308 -128
rect 1298 -137 1308 -133
rect 1312 -133 1317 -128
rect 1312 -137 1322 -133
rect 1336 -133 1342 -128
rect 1331 -137 1342 -133
rect 1346 -133 1350 -128
rect 1346 -137 1355 -133
rect -791 -263 -786 -259
rect -795 -266 -786 -263
rect -783 -263 -774 -259
rect -783 -266 -770 -263
rect -762 -263 -757 -259
rect -766 -266 -757 -263
rect -755 -263 -745 -259
rect -755 -266 -741 -263
rect -733 -263 -726 -259
rect -737 -266 -726 -263
rect -723 -263 -716 -259
rect -723 -266 -712 -263
rect -704 -263 -697 -259
rect -708 -266 -697 -263
rect -694 -263 -687 -259
rect -694 -266 -683 -263
rect -675 -263 -668 -259
rect -679 -266 -668 -263
rect -665 -263 -658 -259
rect -665 -266 -654 -263
rect -646 -263 -638 -259
rect -650 -266 -638 -263
rect -635 -263 -629 -259
rect -635 -266 -625 -263
rect -165 -266 -160 -262
rect -169 -269 -160 -266
rect -157 -266 -148 -262
rect -157 -269 -144 -266
rect -136 -266 -131 -262
rect -140 -269 -131 -266
rect -129 -266 -119 -262
rect -129 -269 -115 -266
rect -107 -266 -100 -262
rect -111 -269 -100 -266
rect -97 -266 -90 -262
rect -97 -269 -86 -266
rect -78 -266 -71 -262
rect -82 -269 -71 -266
rect -68 -266 -61 -262
rect -68 -269 -57 -266
rect -49 -266 -42 -262
rect -53 -269 -42 -266
rect -39 -266 -32 -262
rect -39 -269 -28 -266
rect -20 -266 -12 -262
rect -24 -269 -12 -266
rect -9 -266 -3 -262
rect -9 -269 1 -266
rect 435 -266 440 -262
rect 431 -269 440 -266
rect 443 -266 452 -262
rect 443 -269 456 -266
rect 464 -266 469 -262
rect 460 -269 469 -266
rect 471 -266 481 -262
rect 471 -269 485 -266
rect 493 -266 500 -262
rect 489 -269 500 -266
rect 503 -266 510 -262
rect 503 -269 514 -266
rect 522 -266 529 -262
rect 518 -269 529 -266
rect 532 -266 539 -262
rect 532 -269 543 -266
rect 551 -266 558 -262
rect 547 -269 558 -266
rect 561 -266 568 -262
rect 561 -269 572 -266
rect 580 -266 588 -262
rect 576 -269 588 -266
rect 591 -266 597 -262
rect 1038 -263 1043 -259
rect 1034 -266 1043 -263
rect 1046 -263 1055 -259
rect 1046 -266 1059 -263
rect 1067 -263 1072 -259
rect 1063 -266 1072 -263
rect 1074 -263 1084 -259
rect 1074 -266 1088 -263
rect 1096 -263 1103 -259
rect 1092 -266 1103 -263
rect 1106 -263 1113 -259
rect 1106 -266 1117 -263
rect 1125 -263 1132 -259
rect 1121 -266 1132 -263
rect 1135 -263 1142 -259
rect 1135 -266 1146 -263
rect 1154 -263 1161 -259
rect 1150 -266 1161 -263
rect 1164 -263 1171 -259
rect 1164 -266 1175 -263
rect 1183 -263 1191 -259
rect 1179 -266 1191 -263
rect 1194 -263 1200 -259
rect 1194 -266 1204 -263
rect 591 -269 601 -266
<< pdiffusion >>
rect -830 263 -825 267
rect -834 260 -825 263
rect -822 263 -813 267
rect -822 260 -809 263
rect -801 263 -796 267
rect -805 260 -796 263
rect -794 263 -784 267
rect -794 260 -780 263
rect -772 263 -765 267
rect -776 260 -765 263
rect -762 263 -755 267
rect -762 260 -751 263
rect -743 263 -736 267
rect -747 260 -736 263
rect -733 263 -726 267
rect -733 260 -722 263
rect -714 263 -707 267
rect -718 260 -707 263
rect -704 263 -697 267
rect -704 260 -693 263
rect -685 263 -677 267
rect -689 260 -677 263
rect -674 263 -668 267
rect -674 260 -664 263
rect -612 263 -607 267
rect -616 260 -607 263
rect -604 263 -595 267
rect -604 260 -591 263
rect -583 263 -578 267
rect -587 260 -578 263
rect -576 263 -566 267
rect -576 260 -562 263
rect -554 263 -547 267
rect -558 260 -547 263
rect -544 263 -537 267
rect -544 260 -533 263
rect -525 263 -518 267
rect -529 260 -518 263
rect -515 263 -508 267
rect -515 260 -504 263
rect -496 263 -489 267
rect -500 260 -489 263
rect -486 263 -479 267
rect -486 260 -475 263
rect -467 263 -459 267
rect -471 260 -459 263
rect -456 263 -450 267
rect -456 260 -446 263
rect -379 265 -374 269
rect -383 262 -374 265
rect -371 265 -362 269
rect -371 262 -358 265
rect -350 265 -345 269
rect -354 262 -345 265
rect -343 265 -333 269
rect -343 262 -329 265
rect -321 265 -314 269
rect -325 262 -314 265
rect -311 265 -304 269
rect -311 262 -300 265
rect -292 265 -285 269
rect -296 262 -285 265
rect -282 265 -275 269
rect -282 262 -271 265
rect -263 265 -256 269
rect -267 262 -256 265
rect -253 265 -246 269
rect -253 262 -242 265
rect -234 265 -226 269
rect -238 262 -226 265
rect -223 265 -217 269
rect -223 262 -213 265
rect -119 266 -114 270
rect -123 263 -114 266
rect -111 266 -102 270
rect -111 263 -98 266
rect -90 266 -85 270
rect -94 263 -85 266
rect -83 266 -73 270
rect -83 263 -69 266
rect -61 266 -54 270
rect -65 263 -54 266
rect -51 266 -44 270
rect -51 263 -40 266
rect -32 266 -25 270
rect -36 263 -25 266
rect -22 266 -15 270
rect -22 263 -11 266
rect -3 266 4 270
rect -7 263 4 266
rect 7 266 14 270
rect 7 263 18 266
rect 26 266 34 270
rect 22 263 34 266
rect 37 266 43 270
rect 37 263 47 266
rect -801 65 -796 69
rect -805 62 -796 65
rect -793 65 -784 69
rect -793 62 -780 65
rect -772 65 -767 69
rect -776 62 -767 65
rect -765 65 -755 69
rect -765 62 -751 65
rect -743 65 -736 69
rect -747 62 -736 65
rect -733 65 -726 69
rect -733 62 -722 65
rect -714 65 -707 69
rect -718 62 -707 65
rect -704 65 -697 69
rect -704 62 -693 65
rect -685 65 -678 69
rect -689 62 -678 65
rect -675 65 -668 69
rect -675 62 -664 65
rect -656 65 -648 69
rect -660 62 -648 65
rect -645 65 -639 69
rect -645 62 -635 65
rect -573 64 -569 69
rect -578 60 -569 64
rect -565 64 -559 69
rect -565 60 -554 64
rect -542 64 -537 69
rect -547 60 -537 64
rect -533 64 -528 69
rect -533 60 -523 64
rect -509 64 -503 69
rect -514 60 -503 64
rect -499 64 -495 69
rect -499 60 -490 64
rect -175 62 -170 66
rect -179 59 -170 62
rect -167 62 -158 66
rect -167 59 -154 62
rect -146 62 -141 66
rect -150 59 -141 62
rect -139 62 -129 66
rect -139 59 -125 62
rect -117 62 -110 66
rect -121 59 -110 62
rect -107 62 -100 66
rect -107 59 -96 62
rect -88 62 -81 66
rect -92 59 -81 62
rect -78 62 -71 66
rect -78 59 -67 62
rect -59 62 -52 66
rect -63 59 -52 62
rect -49 62 -42 66
rect -49 59 -38 62
rect -30 62 -22 66
rect -34 59 -22 62
rect -19 62 -13 66
rect -19 59 -9 62
rect 53 61 57 66
rect -398 40 -396 44
rect -394 40 -392 44
rect -380 40 -378 44
rect -376 40 -374 44
rect -361 40 -359 44
rect -357 40 -355 44
rect 48 57 57 61
rect 61 61 67 66
rect 61 57 72 61
rect 84 61 89 66
rect 79 57 89 61
rect 93 61 98 66
rect 93 57 103 61
rect 117 61 123 66
rect 112 57 123 61
rect 127 61 131 66
rect 127 57 136 61
rect 425 62 430 66
rect 421 59 430 62
rect 433 62 442 66
rect 433 59 446 62
rect 454 62 459 66
rect 450 59 459 62
rect 461 62 471 66
rect 461 59 475 62
rect 483 62 490 66
rect 479 59 490 62
rect 493 62 500 66
rect 493 59 504 62
rect 512 62 519 66
rect 508 59 519 62
rect 522 62 529 66
rect 522 59 533 62
rect 541 62 548 66
rect 537 59 548 62
rect 551 62 558 66
rect 551 59 562 62
rect 570 62 578 66
rect 566 59 578 62
rect 581 62 587 66
rect 581 59 591 62
rect 653 61 657 66
rect 228 37 230 41
rect 232 37 234 41
rect 246 37 248 41
rect 250 37 252 41
rect 265 37 267 41
rect 269 37 271 41
rect 648 57 657 61
rect 661 61 667 66
rect 661 57 672 61
rect 684 61 689 66
rect 679 57 689 61
rect 693 61 698 66
rect 693 57 703 61
rect 717 61 723 66
rect 712 57 723 61
rect 727 61 731 66
rect 1028 65 1033 69
rect 1024 62 1033 65
rect 1036 65 1045 69
rect 1036 62 1049 65
rect 1057 65 1062 69
rect 1053 62 1062 65
rect 1064 65 1074 69
rect 1064 62 1078 65
rect 1086 65 1093 69
rect 1082 62 1093 65
rect 1096 65 1103 69
rect 1096 62 1107 65
rect 1115 65 1122 69
rect 1111 62 1122 65
rect 1125 65 1132 69
rect 1125 62 1136 65
rect 1144 65 1151 69
rect 1140 62 1151 65
rect 1154 65 1161 69
rect 1154 62 1165 65
rect 1173 65 1181 69
rect 1169 62 1181 65
rect 1184 65 1190 69
rect 1184 62 1194 65
rect 1256 64 1260 69
rect 727 57 736 61
rect 828 37 830 41
rect 832 37 834 41
rect 846 37 848 41
rect 850 37 852 41
rect 865 37 867 41
rect 869 37 871 41
rect 1251 60 1260 64
rect 1264 64 1270 69
rect 1264 60 1275 64
rect 1287 64 1292 69
rect 1282 60 1292 64
rect 1296 64 1301 69
rect 1296 60 1306 64
rect 1320 64 1326 69
rect 1315 60 1326 64
rect 1330 64 1334 69
rect 1330 60 1339 64
rect 1431 40 1433 44
rect 1435 40 1437 44
rect 1449 40 1451 44
rect 1453 40 1455 44
rect 1468 40 1470 44
rect 1472 40 1474 44
rect -557 -75 -553 -70
rect -562 -79 -553 -75
rect -549 -75 -543 -70
rect -549 -79 -538 -75
rect -526 -75 -521 -70
rect -531 -79 -521 -75
rect -517 -75 -512 -70
rect -517 -79 -507 -75
rect -493 -75 -487 -70
rect -498 -79 -487 -75
rect -483 -75 -479 -70
rect -483 -79 -474 -75
rect 69 -78 73 -73
rect 64 -82 73 -78
rect 77 -78 83 -73
rect 77 -82 88 -78
rect 100 -78 105 -73
rect 95 -82 105 -78
rect 109 -78 114 -73
rect 109 -82 119 -78
rect 133 -78 139 -73
rect 128 -82 139 -78
rect 143 -78 147 -73
rect 143 -82 152 -78
rect 669 -78 673 -73
rect 664 -82 673 -78
rect 677 -78 683 -73
rect 677 -82 688 -78
rect 700 -78 705 -73
rect 695 -82 705 -78
rect 709 -78 714 -73
rect 709 -82 719 -78
rect 733 -78 739 -73
rect 728 -82 739 -78
rect 743 -78 747 -73
rect 743 -82 752 -78
rect 1272 -75 1276 -70
rect 1267 -79 1276 -75
rect 1280 -75 1286 -70
rect 1280 -79 1291 -75
rect 1303 -75 1308 -70
rect 1298 -79 1308 -75
rect 1312 -75 1317 -70
rect 1312 -79 1322 -75
rect 1336 -75 1342 -70
rect 1331 -79 1342 -75
rect 1346 -75 1350 -70
rect 1346 -79 1355 -75
rect -791 -191 -786 -187
rect -795 -194 -786 -191
rect -783 -191 -774 -187
rect -783 -194 -770 -191
rect -762 -191 -757 -187
rect -766 -194 -757 -191
rect -755 -191 -745 -187
rect -755 -194 -741 -191
rect -733 -191 -726 -187
rect -737 -194 -726 -191
rect -723 -191 -716 -187
rect -723 -194 -712 -191
rect -704 -191 -697 -187
rect -708 -194 -697 -191
rect -694 -191 -687 -187
rect -694 -194 -683 -191
rect -675 -191 -668 -187
rect -679 -194 -668 -191
rect -665 -191 -658 -187
rect -665 -194 -654 -191
rect -646 -191 -638 -187
rect -650 -194 -638 -191
rect -635 -191 -629 -187
rect -635 -194 -625 -191
rect -165 -194 -160 -190
rect -169 -197 -160 -194
rect -157 -194 -148 -190
rect -157 -197 -144 -194
rect -136 -194 -131 -190
rect -140 -197 -131 -194
rect -129 -194 -119 -190
rect -129 -197 -115 -194
rect -107 -194 -100 -190
rect -111 -197 -100 -194
rect -97 -194 -90 -190
rect -97 -197 -86 -194
rect -78 -194 -71 -190
rect -82 -197 -71 -194
rect -68 -194 -61 -190
rect -68 -197 -57 -194
rect -49 -194 -42 -190
rect -53 -197 -42 -194
rect -39 -194 -32 -190
rect -39 -197 -28 -194
rect -20 -194 -12 -190
rect -24 -197 -12 -194
rect -9 -194 -3 -190
rect -9 -197 1 -194
rect 435 -194 440 -190
rect 431 -197 440 -194
rect 443 -194 452 -190
rect 443 -197 456 -194
rect 464 -194 469 -190
rect 460 -197 469 -194
rect 471 -194 481 -190
rect 471 -197 485 -194
rect 493 -194 500 -190
rect 489 -197 500 -194
rect 503 -194 510 -190
rect 503 -197 514 -194
rect 522 -194 529 -190
rect 518 -197 529 -194
rect 532 -194 539 -190
rect 532 -197 543 -194
rect 551 -194 558 -190
rect 547 -197 558 -194
rect 561 -194 568 -190
rect 561 -197 572 -194
rect 580 -194 588 -190
rect 576 -197 588 -194
rect 591 -194 597 -190
rect 1038 -191 1043 -187
rect 1034 -194 1043 -191
rect 1046 -191 1055 -187
rect 1046 -194 1059 -191
rect 1067 -191 1072 -187
rect 1063 -194 1072 -191
rect 1074 -191 1084 -187
rect 1074 -194 1088 -191
rect 1096 -191 1103 -187
rect 1092 -194 1103 -191
rect 1106 -191 1113 -187
rect 1106 -194 1117 -191
rect 1125 -191 1132 -187
rect 1121 -194 1132 -191
rect 1135 -191 1142 -187
rect 1135 -194 1146 -191
rect 1154 -191 1161 -187
rect 1150 -194 1161 -191
rect 1164 -191 1171 -187
rect 1164 -194 1175 -191
rect 1183 -191 1191 -187
rect 1179 -194 1191 -191
rect 1194 -191 1200 -187
rect 1194 -194 1204 -191
rect 591 -197 601 -194
<< ndcontact >>
rect -834 191 -830 195
rect -813 191 -809 195
rect -805 191 -801 195
rect -784 191 -780 195
rect -776 191 -772 195
rect -755 191 -751 195
rect -747 191 -743 195
rect -726 191 -722 195
rect -718 191 -714 195
rect -697 191 -693 195
rect -689 191 -685 195
rect -668 191 -664 195
rect -616 191 -612 195
rect -595 191 -591 195
rect -587 191 -583 195
rect -566 191 -562 195
rect -558 191 -554 195
rect -537 191 -533 195
rect -529 191 -525 195
rect -508 191 -504 195
rect -500 191 -496 195
rect -479 191 -475 195
rect -471 191 -467 195
rect -450 191 -446 195
rect -383 193 -379 197
rect -362 193 -358 197
rect -354 193 -350 197
rect -333 193 -329 197
rect -325 193 -321 197
rect -304 193 -300 197
rect -296 193 -292 197
rect -275 193 -271 197
rect -267 193 -263 197
rect -246 193 -242 197
rect -238 193 -234 197
rect -217 193 -213 197
rect -123 194 -119 198
rect -102 194 -98 198
rect -94 194 -90 198
rect -73 194 -69 198
rect -65 194 -61 198
rect -44 194 -40 198
rect -36 194 -32 198
rect -15 194 -11 198
rect -7 194 -3 198
rect 14 194 18 198
rect 22 194 26 198
rect 43 194 47 198
rect -578 6 -573 11
rect -559 6 -554 11
rect -547 6 -542 11
rect -528 6 -523 11
rect -514 6 -509 11
rect -495 6 -490 11
rect -402 -1 -398 3
rect -392 -1 -388 3
rect -384 -1 -380 3
rect -374 -1 -370 3
rect -365 -1 -361 3
rect -355 -1 -351 3
rect -805 -7 -801 -3
rect -784 -7 -780 -3
rect -776 -7 -772 -3
rect -755 -7 -751 -3
rect -747 -7 -743 -3
rect -726 -7 -722 -3
rect -718 -7 -714 -3
rect -697 -7 -693 -3
rect -689 -7 -685 -3
rect -668 -7 -664 -3
rect -660 -7 -656 -3
rect -639 -7 -635 -3
rect 48 3 53 8
rect 67 3 72 8
rect 79 3 84 8
rect 98 3 103 8
rect 112 3 117 8
rect 131 3 136 8
rect 224 -4 228 0
rect 234 -4 238 0
rect 242 -4 246 0
rect 252 -4 256 0
rect 261 -4 265 0
rect 271 -4 275 0
rect -179 -10 -175 -6
rect -158 -10 -154 -6
rect -150 -10 -146 -6
rect -129 -10 -125 -6
rect -121 -10 -117 -6
rect -100 -10 -96 -6
rect -92 -10 -88 -6
rect -71 -10 -67 -6
rect -63 -10 -59 -6
rect -42 -10 -38 -6
rect -34 -10 -30 -6
rect -13 -10 -9 -6
rect 648 3 653 8
rect 667 3 672 8
rect 679 3 684 8
rect 698 3 703 8
rect 712 3 717 8
rect 731 3 736 8
rect 824 -4 828 0
rect 834 -4 838 0
rect 842 -4 846 0
rect 852 -4 856 0
rect 861 -4 865 0
rect 871 -4 875 0
rect 1251 6 1256 11
rect 1270 6 1275 11
rect 1282 6 1287 11
rect 1301 6 1306 11
rect 1315 6 1320 11
rect 1334 6 1339 11
rect 1427 -1 1431 3
rect 1437 -1 1441 3
rect 1445 -1 1449 3
rect 1455 -1 1459 3
rect 1464 -1 1468 3
rect 1474 -1 1478 3
rect 421 -10 425 -6
rect 442 -10 446 -6
rect 450 -10 454 -6
rect 471 -10 475 -6
rect 479 -10 483 -6
rect 500 -10 504 -6
rect 508 -10 512 -6
rect 529 -10 533 -6
rect 537 -10 541 -6
rect 558 -10 562 -6
rect 566 -10 570 -6
rect 587 -10 591 -6
rect 1024 -7 1028 -3
rect 1045 -7 1049 -3
rect 1053 -7 1057 -3
rect 1074 -7 1078 -3
rect 1082 -7 1086 -3
rect 1103 -7 1107 -3
rect 1111 -7 1115 -3
rect 1132 -7 1136 -3
rect 1140 -7 1144 -3
rect 1161 -7 1165 -3
rect 1169 -7 1173 -3
rect 1190 -7 1194 -3
rect -562 -133 -557 -128
rect -543 -133 -538 -128
rect -531 -133 -526 -128
rect -512 -133 -507 -128
rect -498 -133 -493 -128
rect -479 -133 -474 -128
rect 64 -136 69 -131
rect 83 -136 88 -131
rect 95 -136 100 -131
rect 114 -136 119 -131
rect 128 -136 133 -131
rect 147 -136 152 -131
rect 664 -136 669 -131
rect 683 -136 688 -131
rect 695 -136 700 -131
rect 714 -136 719 -131
rect 728 -136 733 -131
rect 747 -136 752 -131
rect 1267 -133 1272 -128
rect 1286 -133 1291 -128
rect 1298 -133 1303 -128
rect 1317 -133 1322 -128
rect 1331 -133 1336 -128
rect 1350 -133 1355 -128
rect -795 -263 -791 -259
rect -774 -263 -770 -259
rect -766 -263 -762 -259
rect -745 -263 -741 -259
rect -737 -263 -733 -259
rect -716 -263 -712 -259
rect -708 -263 -704 -259
rect -687 -263 -683 -259
rect -679 -263 -675 -259
rect -658 -263 -654 -259
rect -650 -263 -646 -259
rect -629 -263 -625 -259
rect -169 -266 -165 -262
rect -148 -266 -144 -262
rect -140 -266 -136 -262
rect -119 -266 -115 -262
rect -111 -266 -107 -262
rect -90 -266 -86 -262
rect -82 -266 -78 -262
rect -61 -266 -57 -262
rect -53 -266 -49 -262
rect -32 -266 -28 -262
rect -24 -266 -20 -262
rect -3 -266 1 -262
rect 431 -266 435 -262
rect 452 -266 456 -262
rect 460 -266 464 -262
rect 481 -266 485 -262
rect 489 -266 493 -262
rect 510 -266 514 -262
rect 518 -266 522 -262
rect 539 -266 543 -262
rect 547 -266 551 -262
rect 568 -266 572 -262
rect 576 -266 580 -262
rect 597 -266 601 -262
rect 1034 -263 1038 -259
rect 1055 -263 1059 -259
rect 1063 -263 1067 -259
rect 1084 -263 1088 -259
rect 1092 -263 1096 -259
rect 1113 -263 1117 -259
rect 1121 -263 1125 -259
rect 1142 -263 1146 -259
rect 1150 -263 1154 -259
rect 1171 -263 1175 -259
rect 1179 -263 1183 -259
rect 1200 -263 1204 -259
<< pdcontact >>
rect -834 263 -830 267
rect -813 263 -809 267
rect -805 263 -801 267
rect -784 263 -780 267
rect -776 263 -772 267
rect -755 263 -751 267
rect -747 263 -743 267
rect -726 263 -722 267
rect -718 263 -714 267
rect -697 263 -693 267
rect -689 263 -685 267
rect -668 263 -664 267
rect -616 263 -612 267
rect -595 263 -591 267
rect -587 263 -583 267
rect -566 263 -562 267
rect -558 263 -554 267
rect -537 263 -533 267
rect -529 263 -525 267
rect -508 263 -504 267
rect -500 263 -496 267
rect -479 263 -475 267
rect -471 263 -467 267
rect -450 263 -446 267
rect -383 265 -379 269
rect -362 265 -358 269
rect -354 265 -350 269
rect -333 265 -329 269
rect -325 265 -321 269
rect -304 265 -300 269
rect -296 265 -292 269
rect -275 265 -271 269
rect -267 265 -263 269
rect -246 265 -242 269
rect -238 265 -234 269
rect -217 265 -213 269
rect -123 266 -119 270
rect -102 266 -98 270
rect -94 266 -90 270
rect -73 266 -69 270
rect -65 266 -61 270
rect -44 266 -40 270
rect -36 266 -32 270
rect -15 266 -11 270
rect -7 266 -3 270
rect 14 266 18 270
rect 22 266 26 270
rect 43 266 47 270
rect -805 65 -801 69
rect -784 65 -780 69
rect -776 65 -772 69
rect -755 65 -751 69
rect -747 65 -743 69
rect -726 65 -722 69
rect -718 65 -714 69
rect -697 65 -693 69
rect -689 65 -685 69
rect -668 65 -664 69
rect -660 65 -656 69
rect -639 65 -635 69
rect -578 64 -573 69
rect -559 64 -554 69
rect -547 64 -542 69
rect -528 64 -523 69
rect -514 64 -509 69
rect -495 64 -490 69
rect -179 62 -175 66
rect -158 62 -154 66
rect -150 62 -146 66
rect -129 62 -125 66
rect -121 62 -117 66
rect -100 62 -96 66
rect -92 62 -88 66
rect -71 62 -67 66
rect -63 62 -59 66
rect -42 62 -38 66
rect -34 62 -30 66
rect -13 62 -9 66
rect 48 61 53 66
rect -402 40 -398 44
rect -392 40 -388 44
rect -384 40 -380 44
rect -374 40 -370 44
rect -365 40 -361 44
rect -355 40 -351 44
rect 67 61 72 66
rect 79 61 84 66
rect 98 61 103 66
rect 112 61 117 66
rect 131 61 136 66
rect 421 62 425 66
rect 442 62 446 66
rect 450 62 454 66
rect 471 62 475 66
rect 479 62 483 66
rect 500 62 504 66
rect 508 62 512 66
rect 529 62 533 66
rect 537 62 541 66
rect 558 62 562 66
rect 566 62 570 66
rect 587 62 591 66
rect 648 61 653 66
rect 224 37 228 41
rect 234 37 238 41
rect 242 37 246 41
rect 252 37 256 41
rect 261 37 265 41
rect 271 37 275 41
rect 667 61 672 66
rect 679 61 684 66
rect 698 61 703 66
rect 712 61 717 66
rect 731 61 736 66
rect 1024 65 1028 69
rect 1045 65 1049 69
rect 1053 65 1057 69
rect 1074 65 1078 69
rect 1082 65 1086 69
rect 1103 65 1107 69
rect 1111 65 1115 69
rect 1132 65 1136 69
rect 1140 65 1144 69
rect 1161 65 1165 69
rect 1169 65 1173 69
rect 1190 65 1194 69
rect 1251 64 1256 69
rect 824 37 828 41
rect 834 37 838 41
rect 842 37 846 41
rect 852 37 856 41
rect 861 37 865 41
rect 871 37 875 41
rect 1270 64 1275 69
rect 1282 64 1287 69
rect 1301 64 1306 69
rect 1315 64 1320 69
rect 1334 64 1339 69
rect 1427 40 1431 44
rect 1437 40 1441 44
rect 1445 40 1449 44
rect 1455 40 1459 44
rect 1464 40 1468 44
rect 1474 40 1478 44
rect -562 -75 -557 -70
rect -543 -75 -538 -70
rect -531 -75 -526 -70
rect -512 -75 -507 -70
rect -498 -75 -493 -70
rect -479 -75 -474 -70
rect 64 -78 69 -73
rect 83 -78 88 -73
rect 95 -78 100 -73
rect 114 -78 119 -73
rect 128 -78 133 -73
rect 147 -78 152 -73
rect 664 -78 669 -73
rect 683 -78 688 -73
rect 695 -78 700 -73
rect 714 -78 719 -73
rect 728 -78 733 -73
rect 747 -78 752 -73
rect 1267 -75 1272 -70
rect 1286 -75 1291 -70
rect 1298 -75 1303 -70
rect 1317 -75 1322 -70
rect 1331 -75 1336 -70
rect 1350 -75 1355 -70
rect -795 -191 -791 -187
rect -774 -191 -770 -187
rect -766 -191 -762 -187
rect -745 -191 -741 -187
rect -737 -191 -733 -187
rect -716 -191 -712 -187
rect -708 -191 -704 -187
rect -687 -191 -683 -187
rect -679 -191 -675 -187
rect -658 -191 -654 -187
rect -650 -191 -646 -187
rect -629 -191 -625 -187
rect -169 -194 -165 -190
rect -148 -194 -144 -190
rect -140 -194 -136 -190
rect -119 -194 -115 -190
rect -111 -194 -107 -190
rect -90 -194 -86 -190
rect -82 -194 -78 -190
rect -61 -194 -57 -190
rect -53 -194 -49 -190
rect -32 -194 -28 -190
rect -24 -194 -20 -190
rect -3 -194 1 -190
rect 431 -194 435 -190
rect 452 -194 456 -190
rect 460 -194 464 -190
rect 481 -194 485 -190
rect 489 -194 493 -190
rect 510 -194 514 -190
rect 518 -194 522 -190
rect 539 -194 543 -190
rect 547 -194 551 -190
rect 568 -194 572 -190
rect 576 -194 580 -190
rect 597 -194 601 -190
rect 1034 -191 1038 -187
rect 1055 -191 1059 -187
rect 1063 -191 1067 -187
rect 1084 -191 1088 -187
rect 1092 -191 1096 -187
rect 1113 -191 1117 -187
rect 1121 -191 1125 -187
rect 1142 -191 1146 -187
rect 1150 -191 1154 -187
rect 1171 -191 1175 -187
rect 1179 -191 1183 -187
rect 1200 -191 1204 -187
<< polysilicon >>
rect -374 275 -311 277
rect -825 273 -762 275
rect -825 267 -822 273
rect -796 267 -794 270
rect -765 267 -762 273
rect -607 273 -544 275
rect -736 267 -733 271
rect -707 267 -704 271
rect -677 267 -674 271
rect -607 267 -604 273
rect -578 267 -576 270
rect -547 267 -544 273
rect -518 267 -515 271
rect -489 267 -486 271
rect -459 267 -456 271
rect -374 269 -371 275
rect -345 269 -343 272
rect -314 269 -311 275
rect -114 276 -51 278
rect -285 269 -282 273
rect -256 269 -253 273
rect -226 269 -223 273
rect -114 270 -111 276
rect -85 270 -83 273
rect -54 270 -51 276
rect -25 270 -22 274
rect 4 270 7 274
rect 34 270 37 274
rect -825 195 -822 260
rect -796 195 -794 260
rect -765 195 -762 260
rect -736 195 -733 260
rect -714 233 -711 238
rect -707 195 -704 260
rect -677 195 -674 260
rect -607 195 -604 260
rect -578 195 -576 260
rect -547 195 -544 260
rect -518 195 -515 260
rect -496 233 -493 238
rect -489 195 -486 260
rect -459 195 -456 260
rect -374 197 -371 262
rect -345 197 -343 262
rect -314 197 -311 262
rect -285 197 -282 262
rect -263 235 -260 240
rect -256 197 -253 262
rect -226 197 -223 262
rect -114 198 -111 263
rect -85 198 -83 263
rect -54 198 -51 263
rect -25 198 -22 263
rect -3 236 0 241
rect 4 198 7 263
rect 34 198 37 263
rect -825 183 -822 188
rect -796 176 -794 188
rect -765 185 -762 188
rect -736 176 -733 188
rect -707 183 -704 188
rect -677 183 -674 188
rect -607 183 -604 188
rect -796 174 -733 176
rect -578 176 -576 188
rect -547 185 -544 188
rect -518 176 -515 188
rect -489 183 -486 188
rect -459 183 -456 188
rect -374 185 -371 190
rect -578 173 -515 176
rect -345 178 -343 190
rect -314 187 -311 190
rect -285 178 -282 190
rect -256 185 -253 190
rect -226 185 -223 190
rect -114 186 -111 191
rect -345 175 -282 178
rect -85 179 -83 191
rect -54 188 -51 191
rect -25 179 -22 191
rect 4 186 7 191
rect 34 186 37 191
rect -85 176 -22 179
rect -796 75 -733 77
rect 1033 75 1096 77
rect -796 69 -793 75
rect -767 69 -765 72
rect -736 69 -733 75
rect -707 69 -704 73
rect -678 69 -675 73
rect -648 69 -645 73
rect -569 69 -565 75
rect -537 69 -533 73
rect -503 69 -499 73
rect -170 72 -107 74
rect 430 72 493 74
rect -796 -3 -793 62
rect -767 -3 -765 62
rect -736 -3 -733 62
rect -707 -3 -704 62
rect -685 35 -682 40
rect -678 -3 -675 62
rect -648 -3 -645 62
rect -170 66 -167 72
rect -141 66 -139 69
rect -110 66 -107 72
rect -81 66 -78 70
rect -52 66 -49 70
rect -22 66 -19 70
rect 57 66 61 72
rect 89 66 93 70
rect 123 66 127 70
rect 430 66 433 72
rect 459 66 461 69
rect 490 66 493 72
rect 519 66 522 70
rect 548 66 551 70
rect 578 66 581 70
rect 657 66 661 72
rect 689 66 693 70
rect 723 66 727 70
rect 1033 69 1036 75
rect 1062 69 1064 72
rect 1093 69 1096 75
rect 1122 69 1125 73
rect 1151 69 1154 73
rect 1181 69 1184 73
rect 1260 69 1264 75
rect 1292 69 1296 73
rect 1326 69 1330 73
rect -569 26 -565 60
rect -568 21 -565 26
rect -569 11 -565 21
rect -537 11 -533 60
rect -503 11 -499 60
rect -396 44 -394 47
rect -378 44 -376 47
rect -359 44 -357 47
rect -396 17 -394 40
rect -378 19 -376 40
rect -359 20 -357 40
rect -395 13 -394 17
rect -377 15 -376 19
rect -358 16 -357 20
rect -396 3 -394 13
rect -378 3 -376 15
rect -359 3 -357 16
rect -569 -1 -565 2
rect -537 -1 -533 2
rect -503 -1 -499 2
rect -396 -4 -394 -1
rect -378 -4 -376 -1
rect -359 -4 -357 -1
rect -170 -6 -167 59
rect -141 -6 -139 59
rect -110 -6 -107 59
rect -81 -6 -78 59
rect -59 32 -56 37
rect -52 -6 -49 59
rect -22 -6 -19 59
rect 57 23 61 57
rect 58 18 61 23
rect 57 8 61 18
rect 89 8 93 57
rect 123 8 127 57
rect 230 41 232 44
rect 248 41 250 44
rect 267 41 269 44
rect 230 14 232 37
rect 248 16 250 37
rect 267 17 269 37
rect 231 10 232 14
rect 249 12 250 16
rect 268 13 269 17
rect 230 0 232 10
rect 248 0 250 12
rect 267 0 269 13
rect 57 -4 61 -1
rect 89 -4 93 -1
rect 123 -4 127 -1
rect -796 -15 -793 -10
rect -767 -22 -765 -10
rect -736 -13 -733 -10
rect -707 -22 -704 -10
rect -678 -15 -675 -10
rect -648 -15 -645 -10
rect 230 -7 232 -4
rect 248 -7 250 -4
rect 267 -7 269 -4
rect 430 -6 433 59
rect 459 -6 461 59
rect 490 -6 493 59
rect 519 -6 522 59
rect 541 32 544 37
rect 548 -6 551 59
rect 578 -6 581 59
rect 657 23 661 57
rect 658 18 661 23
rect 657 8 661 18
rect 689 8 693 57
rect 723 8 727 57
rect 830 41 832 44
rect 848 41 850 44
rect 867 41 869 44
rect 830 14 832 37
rect 848 16 850 37
rect 867 17 869 37
rect 831 10 832 14
rect 849 12 850 16
rect 868 13 869 17
rect 830 0 832 10
rect 848 0 850 12
rect 867 0 869 13
rect 657 -4 661 -1
rect 689 -4 693 -1
rect 723 -4 727 -1
rect 1033 -3 1036 62
rect 1062 -3 1064 62
rect 1093 -3 1096 62
rect 1122 -3 1125 62
rect 1144 35 1147 40
rect 1151 -3 1154 62
rect 1181 -3 1184 62
rect 1260 26 1264 60
rect 1261 21 1264 26
rect 1260 11 1264 21
rect 1292 11 1296 60
rect 1326 11 1330 60
rect 1433 44 1435 47
rect 1451 44 1453 47
rect 1470 44 1472 47
rect 1433 17 1435 40
rect 1451 19 1453 40
rect 1470 20 1472 40
rect 1434 13 1435 17
rect 1452 15 1453 19
rect 1471 16 1472 20
rect 1433 3 1435 13
rect 1451 3 1453 15
rect 1470 3 1472 16
rect 1260 -1 1264 2
rect 1292 -1 1296 2
rect 1326 -1 1330 2
rect 830 -7 832 -4
rect 848 -7 850 -4
rect 867 -7 869 -4
rect 1433 -4 1435 -1
rect 1451 -4 1453 -1
rect 1470 -4 1472 -1
rect -170 -18 -167 -13
rect -767 -25 -704 -22
rect -141 -25 -139 -13
rect -110 -16 -107 -13
rect -81 -25 -78 -13
rect -52 -18 -49 -13
rect -22 -18 -19 -13
rect 430 -18 433 -13
rect -141 -28 -78 -25
rect 459 -25 461 -13
rect 490 -16 493 -13
rect 519 -25 522 -13
rect 548 -18 551 -13
rect 578 -18 581 -13
rect 1033 -15 1036 -10
rect 1062 -22 1064 -10
rect 1093 -13 1096 -10
rect 1122 -22 1125 -10
rect 1151 -15 1154 -10
rect 1181 -15 1184 -10
rect 1062 -25 1125 -22
rect 459 -28 522 -25
rect -553 -70 -549 -64
rect -521 -70 -517 -66
rect -487 -70 -483 -66
rect 73 -73 77 -67
rect 105 -73 109 -69
rect 139 -73 143 -69
rect 673 -73 677 -67
rect 705 -73 709 -69
rect 739 -73 743 -69
rect 1276 -70 1280 -64
rect 1308 -70 1312 -66
rect 1342 -70 1346 -66
rect -553 -113 -549 -79
rect -552 -118 -549 -113
rect -553 -128 -549 -118
rect -521 -128 -517 -79
rect -487 -128 -483 -79
rect 73 -116 77 -82
rect 74 -121 77 -116
rect 73 -131 77 -121
rect 105 -131 109 -82
rect 139 -131 143 -82
rect 673 -116 677 -82
rect 674 -121 677 -116
rect 673 -131 677 -121
rect 705 -131 709 -82
rect 739 -131 743 -82
rect 1276 -113 1280 -79
rect 1277 -118 1280 -113
rect 1276 -128 1280 -118
rect 1308 -128 1312 -79
rect 1342 -128 1346 -79
rect -553 -140 -549 -137
rect -521 -140 -517 -137
rect -487 -140 -483 -137
rect 1276 -140 1280 -137
rect 1308 -140 1312 -137
rect 1342 -140 1346 -137
rect 73 -143 77 -140
rect 105 -143 109 -140
rect 139 -143 143 -140
rect 673 -143 677 -140
rect 705 -143 709 -140
rect 739 -143 743 -140
rect -786 -181 -723 -179
rect -786 -187 -783 -181
rect -757 -187 -755 -184
rect -726 -187 -723 -181
rect 1043 -181 1106 -179
rect -697 -187 -694 -183
rect -668 -187 -665 -183
rect -638 -187 -635 -183
rect -160 -184 -97 -182
rect -160 -190 -157 -184
rect -131 -190 -129 -187
rect -100 -190 -97 -184
rect 440 -184 503 -182
rect -71 -190 -68 -186
rect -42 -190 -39 -186
rect -12 -190 -9 -186
rect 440 -190 443 -184
rect 469 -190 471 -187
rect 500 -190 503 -184
rect 529 -190 532 -186
rect 558 -190 561 -186
rect 588 -190 591 -186
rect 1043 -187 1046 -181
rect 1072 -187 1074 -184
rect 1103 -187 1106 -181
rect 1132 -187 1135 -183
rect 1161 -187 1164 -183
rect 1191 -187 1194 -183
rect -786 -259 -783 -194
rect -757 -259 -755 -194
rect -726 -259 -723 -194
rect -697 -259 -694 -194
rect -675 -221 -672 -216
rect -668 -259 -665 -194
rect -638 -259 -635 -194
rect -160 -262 -157 -197
rect -131 -262 -129 -197
rect -100 -262 -97 -197
rect -71 -262 -68 -197
rect -49 -224 -46 -219
rect -42 -262 -39 -197
rect -12 -262 -9 -197
rect 440 -262 443 -197
rect 469 -262 471 -197
rect 500 -262 503 -197
rect 529 -262 532 -197
rect 551 -224 554 -219
rect 558 -262 561 -197
rect 588 -262 591 -197
rect 1043 -259 1046 -194
rect 1072 -259 1074 -194
rect 1103 -259 1106 -194
rect 1132 -259 1135 -194
rect 1154 -221 1157 -216
rect 1161 -259 1164 -194
rect 1191 -259 1194 -194
rect -786 -271 -783 -266
rect -757 -278 -755 -266
rect -726 -269 -723 -266
rect -697 -278 -694 -266
rect -668 -271 -665 -266
rect -638 -271 -635 -266
rect -160 -274 -157 -269
rect -757 -281 -694 -278
rect -131 -281 -129 -269
rect -100 -272 -97 -269
rect -71 -281 -68 -269
rect -42 -274 -39 -269
rect -12 -274 -9 -269
rect 440 -274 443 -269
rect -131 -284 -68 -281
rect 469 -281 471 -269
rect 500 -272 503 -269
rect 529 -281 532 -269
rect 558 -274 561 -269
rect 588 -274 591 -269
rect 1043 -271 1046 -266
rect 1072 -278 1074 -266
rect 1103 -269 1106 -266
rect 1132 -278 1135 -266
rect 1161 -271 1164 -266
rect 1191 -271 1194 -266
rect 1072 -281 1135 -278
rect 469 -284 532 -281
<< polycontact >>
rect -830 224 -825 229
rect -801 223 -796 228
rect -711 233 -707 238
rect -682 206 -677 212
rect -612 224 -607 229
rect -583 223 -578 228
rect -493 233 -489 238
rect -464 206 -459 212
rect -379 226 -374 231
rect -350 225 -345 230
rect -260 235 -256 240
rect -231 208 -226 214
rect -119 227 -114 232
rect -90 226 -85 231
rect 0 236 4 241
rect 29 209 34 215
rect -801 26 -796 31
rect -772 25 -767 30
rect -682 35 -678 40
rect -653 8 -648 14
rect -572 21 -568 26
rect -541 21 -537 26
rect -509 34 -503 40
rect -175 23 -170 28
rect -399 13 -395 17
rect -381 15 -377 19
rect -362 16 -358 20
rect -146 22 -141 27
rect -56 32 -52 37
rect -27 5 -22 11
rect 54 18 58 23
rect 85 18 89 23
rect 117 31 123 37
rect 425 23 430 28
rect 227 10 231 14
rect 245 12 249 16
rect 264 13 268 17
rect 454 22 459 27
rect 544 32 548 37
rect 573 5 578 11
rect 654 18 658 23
rect 685 18 689 23
rect 717 31 723 37
rect 1028 26 1033 31
rect 827 10 831 14
rect 845 12 849 16
rect 864 13 868 17
rect 1057 25 1062 30
rect 1147 35 1151 40
rect 1176 8 1181 14
rect 1257 21 1261 26
rect 1288 21 1292 26
rect 1320 34 1326 40
rect 1430 13 1434 17
rect 1448 15 1452 19
rect 1467 16 1471 20
rect -556 -118 -552 -113
rect -525 -118 -521 -113
rect -493 -105 -487 -99
rect 70 -121 74 -116
rect 101 -121 105 -116
rect 133 -108 139 -102
rect 670 -121 674 -116
rect 701 -121 705 -116
rect 733 -108 739 -102
rect 1273 -118 1277 -113
rect 1304 -118 1308 -113
rect 1336 -105 1342 -99
rect -791 -230 -786 -225
rect -762 -231 -757 -226
rect -672 -221 -668 -216
rect -643 -248 -638 -242
rect -165 -233 -160 -228
rect -136 -234 -131 -229
rect -46 -224 -42 -219
rect -17 -251 -12 -245
rect 435 -233 440 -228
rect 464 -234 469 -229
rect 554 -224 558 -219
rect 583 -251 588 -245
rect 1038 -230 1043 -225
rect 1067 -231 1072 -226
rect 1157 -221 1161 -216
rect 1186 -248 1191 -242
<< metal1 >>
rect -389 294 59 295
rect -440 293 59 294
rect -869 289 59 293
rect -869 288 -201 289
rect -869 287 -365 288
rect -869 277 -862 287
rect -840 286 -434 287
rect -868 94 -862 277
rect -834 267 -830 286
rect -805 267 -801 286
rect -776 267 -772 286
rect -747 267 -743 286
rect -726 272 -685 276
rect -726 267 -722 272
rect -718 267 -714 272
rect -689 267 -685 272
rect -616 267 -612 286
rect -587 267 -583 286
rect -558 267 -554 286
rect -529 267 -525 286
rect -508 272 -467 276
rect -508 267 -504 272
rect -500 267 -496 272
rect -471 267 -467 272
rect -383 269 -379 287
rect -354 269 -350 288
rect -325 269 -321 288
rect -296 269 -292 288
rect -275 274 -234 278
rect -275 269 -271 274
rect -267 269 -263 274
rect -238 269 -234 274
rect -123 270 -119 289
rect -94 270 -90 289
rect -65 270 -61 289
rect -36 270 -32 289
rect -15 275 26 279
rect -15 270 -11 275
rect -7 270 -3 275
rect 22 270 26 275
rect -833 224 -830 229
rect -813 195 -809 263
rect -806 223 -801 228
rect -784 212 -780 263
rect -755 256 -751 263
rect -726 256 -722 263
rect -755 253 -722 256
rect -697 256 -693 263
rect -668 256 -664 263
rect -697 253 -664 256
rect -719 234 -711 238
rect -714 233 -711 234
rect -668 230 -664 253
rect -668 229 -653 230
rect -668 220 -662 229
rect -613 224 -612 229
rect -784 207 -682 212
rect -784 195 -780 207
rect -686 206 -682 207
rect -668 203 -664 220
rect -726 195 -722 196
rect -668 195 -664 198
rect -595 195 -591 263
rect -588 223 -583 228
rect -566 212 -562 263
rect -537 256 -533 263
rect -508 256 -504 263
rect -537 253 -504 256
rect -479 256 -475 263
rect -450 256 -446 263
rect -479 253 -446 256
rect -501 234 -493 238
rect -496 233 -493 234
rect -566 207 -464 212
rect -566 195 -562 207
rect -468 206 -464 207
rect -450 203 -446 253
rect -382 226 -379 231
rect -508 195 -504 196
rect -450 195 -446 198
rect -362 197 -358 265
rect -355 225 -350 230
rect -333 214 -329 265
rect -304 258 -300 265
rect -275 258 -271 265
rect -304 255 -271 258
rect -246 258 -242 265
rect -217 258 -213 265
rect -246 255 -213 258
rect -268 236 -260 240
rect -263 235 -260 236
rect -217 232 -213 255
rect -217 222 -181 232
rect -122 227 -119 232
rect -333 209 -231 214
rect -333 197 -329 209
rect -235 208 -231 209
rect -217 205 -213 222
rect -275 197 -271 198
rect -217 197 -213 200
rect -102 198 -98 266
rect -95 226 -90 231
rect -73 215 -69 266
rect -44 259 -40 266
rect -15 259 -11 266
rect -44 256 -11 259
rect 14 259 18 266
rect 43 259 47 266
rect 14 256 47 259
rect -8 237 0 241
rect -3 236 0 237
rect 43 233 47 256
rect 43 232 51 233
rect 43 224 92 232
rect 43 223 51 224
rect -73 210 29 215
rect -73 198 -69 210
rect 25 209 29 210
rect 43 206 47 223
rect -15 198 -11 199
rect 43 198 47 201
rect -751 191 -747 195
rect -693 191 -689 195
rect -533 191 -529 195
rect -475 191 -471 195
rect -300 193 -296 197
rect -242 193 -238 197
rect -40 194 -36 198
rect 18 194 22 198
rect -834 187 -830 191
rect -805 187 -801 191
rect -776 187 -772 191
rect -718 187 -714 191
rect -616 187 -612 191
rect -587 187 -583 191
rect -558 187 -554 191
rect -500 187 -496 191
rect -383 189 -379 193
rect -354 189 -350 193
rect -325 189 -321 193
rect -267 189 -263 193
rect -386 188 -198 189
rect -437 187 -128 188
rect -123 187 -119 194
rect -94 190 -90 194
rect -65 190 -61 194
rect -7 190 -3 194
rect -116 189 62 190
rect -116 187 1609 189
rect -837 183 1609 187
rect -837 182 -107 183
rect 54 182 1609 183
rect -837 181 -382 182
rect -837 180 -431 181
rect -868 88 -598 94
rect -141 91 -137 92
rect -242 88 28 91
rect -868 87 -795 88
rect -868 -154 -854 87
rect -805 69 -801 87
rect -776 69 -772 88
rect -747 69 -743 88
rect -718 69 -714 88
rect -603 85 -598 88
rect -353 85 28 88
rect -603 84 -169 85
rect -603 79 -228 84
rect -603 78 -330 79
rect -697 74 -656 78
rect -697 69 -693 74
rect -689 69 -685 74
rect -660 69 -656 74
rect -578 69 -573 78
rect -547 69 -542 78
rect -514 69 -509 78
rect -784 41 -780 65
rect -784 37 -764 41
rect -803 26 -801 31
rect -784 -3 -780 37
rect -755 14 -751 65
rect -726 58 -722 65
rect -697 58 -693 65
rect -726 55 -693 58
rect -668 58 -664 65
rect -639 58 -635 65
rect -668 55 -635 58
rect -690 36 -682 40
rect -685 35 -682 36
rect -639 32 -635 55
rect -559 40 -554 64
rect -528 40 -523 64
rect -559 34 -509 40
rect -639 29 -631 32
rect -639 24 -597 29
rect -639 22 -631 24
rect -755 9 -653 14
rect -755 -3 -751 9
rect -657 8 -653 9
rect -639 5 -635 22
rect -697 -3 -693 -2
rect -639 -3 -635 0
rect -722 -7 -718 -3
rect -664 -7 -660 -3
rect -805 -11 -801 -7
rect -776 -11 -772 -7
rect -747 -10 -743 -7
rect -749 -11 -743 -10
rect -689 -11 -685 -7
rect -833 -18 -627 -11
rect -833 -267 -821 -18
rect -604 -113 -597 24
rect -573 21 -572 26
rect -542 21 -541 26
rect -528 11 -523 34
rect -495 11 -490 64
rect -336 55 -330 78
rect -416 50 -330 55
rect -402 44 -398 50
rect -365 44 -361 50
rect -388 40 -384 44
rect -374 20 -370 40
rect -355 26 -351 40
rect -554 6 -547 11
rect -421 13 -399 17
rect -382 15 -381 19
rect -374 16 -362 20
rect -355 19 -352 26
rect -421 12 -400 13
rect -578 2 -573 6
rect -514 2 -509 6
rect -584 1 -483 2
rect -577 -5 -483 1
rect -569 -61 -440 -54
rect -562 -70 -557 -61
rect -531 -70 -526 -61
rect -498 -70 -493 -61
rect -543 -99 -538 -75
rect -512 -99 -507 -75
rect -543 -105 -493 -99
rect -479 -102 -474 -75
rect -421 -102 -414 12
rect -374 11 -370 16
rect -392 8 -370 11
rect -392 3 -388 8
rect -374 3 -370 8
rect -355 3 -351 19
rect -402 -4 -398 -1
rect -384 -4 -380 -1
rect -365 -4 -361 -1
rect -406 -5 -342 -4
rect -397 -7 -342 -5
rect -337 -54 -330 50
rect -374 -61 -330 -54
rect -604 -118 -556 -113
rect -528 -118 -525 -113
rect -793 -167 -613 -161
rect -801 -168 -613 -167
rect -795 -187 -791 -168
rect -766 -187 -762 -168
rect -737 -187 -733 -168
rect -708 -187 -704 -168
rect -687 -182 -646 -178
rect -687 -187 -683 -182
rect -679 -187 -675 -182
rect -650 -187 -646 -182
rect -794 -230 -791 -225
rect -774 -259 -770 -191
rect -745 -242 -741 -191
rect -716 -198 -712 -191
rect -687 -198 -683 -191
rect -716 -201 -683 -198
rect -658 -198 -654 -191
rect -629 -198 -625 -191
rect -658 -201 -625 -198
rect -680 -220 -672 -216
rect -675 -221 -672 -220
rect -629 -224 -625 -201
rect -629 -234 -621 -224
rect -745 -247 -643 -242
rect -745 -259 -741 -247
rect -647 -248 -643 -247
rect -629 -251 -625 -234
rect -687 -259 -683 -258
rect -629 -259 -625 -256
rect -712 -263 -708 -259
rect -654 -263 -650 -259
rect -795 -267 -791 -263
rect -766 -267 -762 -263
rect -737 -267 -733 -263
rect -679 -267 -675 -263
rect -833 -274 -610 -267
rect -833 -332 -821 -274
rect -604 -295 -597 -118
rect -512 -128 -507 -105
rect -479 -107 -414 -102
rect -479 -128 -474 -107
rect -538 -133 -531 -128
rect -562 -137 -557 -133
rect -498 -137 -493 -133
rect -760 -302 -597 -295
rect -568 -144 -461 -137
rect -568 -332 -554 -144
rect -242 -157 -228 79
rect -179 66 -175 84
rect -150 66 -146 85
rect -121 66 -117 85
rect -92 66 -88 85
rect 23 82 28 85
rect 358 85 628 91
rect 358 84 431 85
rect 358 83 372 84
rect 291 82 372 83
rect 23 75 372 82
rect -71 71 -30 75
rect -71 66 -67 71
rect -63 66 -59 71
rect -34 66 -30 71
rect 48 66 53 75
rect 79 66 84 75
rect 112 66 117 75
rect -158 38 -154 62
rect -158 34 -138 38
rect -177 23 -175 28
rect -158 -6 -154 34
rect -129 11 -125 62
rect -100 55 -96 62
rect -71 55 -67 62
rect -100 52 -67 55
rect -42 55 -38 62
rect -13 55 -9 62
rect -42 52 -9 55
rect -64 33 -56 37
rect -59 32 -56 33
rect -13 29 -9 52
rect 67 37 72 61
rect 98 37 103 61
rect 67 31 117 37
rect -13 26 -5 29
rect -13 21 29 26
rect -13 19 -5 21
rect -129 6 -27 11
rect -129 -6 -125 6
rect -31 5 -27 6
rect -13 2 -9 19
rect -71 -6 -67 -5
rect -13 -6 -9 -3
rect -96 -10 -92 -6
rect -38 -10 -34 -6
rect -179 -14 -175 -10
rect -150 -14 -146 -10
rect -121 -14 -117 -10
rect -63 -14 -59 -10
rect -207 -21 -1 -14
rect -833 -335 -554 -332
rect -207 -270 -195 -21
rect 22 -116 29 21
rect 53 18 54 23
rect 84 18 85 23
rect 98 8 103 31
rect 131 8 136 61
rect 290 52 296 75
rect 210 47 296 52
rect 224 41 228 47
rect 261 41 265 47
rect 238 37 242 41
rect 252 17 256 37
rect 271 20 275 37
rect 72 3 79 8
rect 205 10 227 14
rect 244 12 245 16
rect 252 13 264 17
rect 271 16 278 20
rect 205 9 226 10
rect 48 -1 53 3
rect 112 -1 117 3
rect 42 -2 143 -1
rect 49 -8 143 -2
rect 57 -64 186 -57
rect 64 -73 69 -64
rect 95 -73 100 -64
rect 128 -73 133 -64
rect 83 -102 88 -78
rect 114 -102 119 -78
rect 83 -108 133 -102
rect 147 -105 152 -78
rect 205 -105 212 9
rect 252 8 256 13
rect 234 5 256 8
rect 234 0 238 5
rect 252 0 256 5
rect 271 0 275 16
rect 224 -7 228 -4
rect 242 -7 246 -4
rect 261 -7 265 -4
rect 220 -8 284 -7
rect 229 -10 284 -8
rect 289 -57 296 47
rect 252 -64 296 -57
rect 22 -121 70 -116
rect 98 -121 101 -116
rect -167 -170 13 -164
rect -175 -171 13 -170
rect -169 -190 -165 -171
rect -140 -190 -136 -171
rect -111 -190 -107 -171
rect -82 -190 -78 -171
rect -61 -185 -20 -181
rect -61 -190 -57 -185
rect -53 -190 -49 -185
rect -24 -190 -20 -185
rect -168 -233 -165 -228
rect -148 -262 -144 -194
rect -119 -245 -115 -194
rect -90 -201 -86 -194
rect -61 -201 -57 -194
rect -90 -204 -57 -201
rect -32 -201 -28 -194
rect -3 -201 1 -194
rect -32 -204 1 -201
rect -54 -223 -46 -219
rect -49 -224 -46 -223
rect -3 -227 1 -204
rect -3 -237 5 -227
rect -119 -250 -17 -245
rect -119 -262 -115 -250
rect -21 -251 -17 -250
rect -3 -254 1 -237
rect -61 -262 -57 -261
rect -3 -262 1 -259
rect -86 -266 -82 -262
rect -28 -266 -24 -262
rect -169 -270 -165 -266
rect -140 -270 -136 -266
rect -111 -270 -107 -266
rect -53 -270 -49 -266
rect -207 -277 16 -270
rect -207 -335 -195 -277
rect 22 -298 29 -121
rect 114 -131 119 -108
rect 147 -110 212 -105
rect 147 -131 152 -110
rect 88 -136 95 -131
rect 64 -140 69 -136
rect 128 -140 133 -136
rect -134 -305 29 -298
rect 58 -147 165 -140
rect 58 -335 72 -147
rect 358 -157 372 75
rect 421 66 425 84
rect 450 66 454 85
rect 458 84 462 85
rect 479 66 483 85
rect 508 66 512 85
rect 623 82 628 85
rect 961 88 1231 94
rect 961 87 1034 88
rect 623 77 896 82
rect 961 77 975 87
rect 623 75 975 77
rect 529 71 570 75
rect 529 66 533 71
rect 537 66 541 71
rect 566 66 570 71
rect 648 66 653 75
rect 679 66 684 75
rect 712 66 717 75
rect 890 69 975 75
rect 442 38 446 62
rect 442 34 462 38
rect 423 23 425 28
rect 442 -6 446 34
rect 471 11 475 62
rect 500 55 504 62
rect 529 55 533 62
rect 500 52 533 55
rect 558 55 562 62
rect 587 55 591 62
rect 558 52 591 55
rect 536 33 544 37
rect 541 32 544 33
rect 587 29 591 52
rect 667 37 672 61
rect 698 37 703 61
rect 667 31 717 37
rect 587 26 595 29
rect 587 21 629 26
rect 587 19 595 21
rect 471 6 573 11
rect 471 -6 475 6
rect 569 5 573 6
rect 587 2 591 19
rect 529 -6 533 -5
rect 587 -6 591 -3
rect 504 -10 508 -6
rect 562 -10 566 -6
rect 421 -14 425 -10
rect 450 -14 454 -10
rect 479 -14 483 -10
rect 537 -14 541 -10
rect 393 -21 599 -14
rect -833 -339 72 -335
rect 393 -270 405 -21
rect 622 -116 629 21
rect 653 18 654 23
rect 684 18 685 23
rect 698 8 703 31
rect 731 8 736 61
rect 890 52 896 69
rect 810 47 896 52
rect 824 41 828 47
rect 861 41 865 47
rect 838 37 842 41
rect 852 17 856 37
rect 871 20 875 37
rect 672 3 679 8
rect 805 10 827 14
rect 844 12 845 16
rect 852 13 864 17
rect 871 16 878 20
rect 805 9 826 10
rect 648 -1 653 3
rect 712 -1 717 3
rect 642 -2 743 -1
rect 649 -8 743 -2
rect 657 -64 786 -57
rect 664 -73 669 -64
rect 695 -73 700 -64
rect 728 -73 733 -64
rect 683 -102 688 -78
rect 714 -102 719 -78
rect 683 -108 733 -102
rect 747 -105 752 -78
rect 805 -105 812 9
rect 852 8 856 13
rect 834 5 856 8
rect 834 0 838 5
rect 852 0 856 5
rect 871 0 875 16
rect 824 -7 828 -4
rect 842 -7 846 -4
rect 861 -7 865 -4
rect 820 -8 884 -7
rect 829 -10 884 -8
rect 889 -57 896 47
rect 852 -64 896 -57
rect 622 -121 670 -116
rect 698 -121 701 -116
rect 433 -170 613 -164
rect 425 -171 613 -170
rect 431 -190 435 -171
rect 460 -190 464 -171
rect 489 -190 493 -171
rect 518 -190 522 -171
rect 539 -185 580 -181
rect 539 -190 543 -185
rect 547 -190 551 -185
rect 576 -190 580 -185
rect 433 -233 435 -228
rect 452 -262 456 -194
rect 481 -245 485 -194
rect 510 -201 514 -194
rect 539 -201 543 -194
rect 510 -204 543 -201
rect 568 -201 572 -194
rect 597 -201 601 -194
rect 568 -204 601 -201
rect 546 -223 554 -219
rect 551 -224 554 -223
rect 597 -227 601 -204
rect 597 -237 605 -227
rect 481 -250 583 -245
rect 481 -262 485 -250
rect 579 -251 583 -250
rect 597 -254 601 -237
rect 539 -262 543 -261
rect 597 -262 601 -259
rect 514 -266 518 -262
rect 572 -266 576 -262
rect 431 -270 435 -266
rect 460 -270 464 -266
rect 489 -270 493 -266
rect 547 -270 551 -266
rect 393 -277 616 -270
rect 393 -335 405 -277
rect 622 -298 629 -121
rect 714 -131 719 -108
rect 747 -110 812 -105
rect 747 -131 752 -110
rect 688 -136 695 -131
rect 664 -140 669 -136
rect 728 -140 733 -136
rect 466 -305 629 -298
rect 658 -147 765 -140
rect 658 -335 672 -147
rect 961 -154 975 69
rect 1024 69 1028 87
rect 1053 69 1057 88
rect 1082 69 1086 88
rect 1111 69 1115 88
rect 1226 85 1231 88
rect 1226 78 1499 85
rect 1132 74 1173 78
rect 1132 69 1136 74
rect 1140 69 1144 74
rect 1169 69 1173 74
rect 1251 69 1256 78
rect 1282 69 1287 78
rect 1315 69 1320 78
rect 1045 41 1049 65
rect 1045 37 1065 41
rect 1026 26 1028 31
rect 1045 -3 1049 37
rect 1074 14 1078 65
rect 1103 58 1107 65
rect 1132 58 1136 65
rect 1103 55 1136 58
rect 1161 58 1165 65
rect 1190 58 1194 65
rect 1161 55 1194 58
rect 1139 36 1147 40
rect 1144 35 1147 36
rect 1190 32 1194 55
rect 1270 40 1275 64
rect 1301 40 1306 64
rect 1270 34 1320 40
rect 1190 29 1198 32
rect 1190 24 1232 29
rect 1190 22 1198 24
rect 1074 9 1176 14
rect 1074 -3 1078 9
rect 1172 8 1176 9
rect 1190 5 1194 22
rect 1132 -3 1136 -2
rect 1190 -3 1194 0
rect 1107 -7 1111 -3
rect 1165 -7 1169 -3
rect 1024 -11 1028 -7
rect 1053 -11 1057 -7
rect 1082 -9 1086 -7
rect 1081 -11 1086 -9
rect 1140 -11 1144 -7
rect 996 -18 1202 -11
rect 393 -336 672 -335
rect 996 -267 1008 -18
rect 1225 -113 1232 24
rect 1256 21 1257 26
rect 1287 21 1288 26
rect 1301 11 1306 34
rect 1334 11 1339 64
rect 1493 55 1499 78
rect 1413 50 1499 55
rect 1427 44 1431 50
rect 1464 44 1468 50
rect 1441 40 1445 44
rect 1455 20 1459 40
rect 1474 23 1478 40
rect 1275 6 1282 11
rect 1408 13 1430 17
rect 1447 15 1448 19
rect 1455 16 1467 20
rect 1474 19 1483 23
rect 1408 12 1429 13
rect 1251 2 1256 6
rect 1315 2 1320 6
rect 1245 1 1346 2
rect 1252 -5 1346 1
rect 1260 -61 1389 -54
rect 1267 -70 1272 -61
rect 1298 -70 1303 -61
rect 1331 -70 1336 -61
rect 1286 -99 1291 -75
rect 1317 -99 1322 -75
rect 1286 -105 1336 -99
rect 1350 -102 1355 -75
rect 1408 -102 1415 12
rect 1455 11 1459 16
rect 1437 8 1459 11
rect 1437 3 1441 8
rect 1455 3 1459 8
rect 1474 3 1478 19
rect 1427 -4 1431 -1
rect 1445 -4 1449 -1
rect 1464 -4 1468 -1
rect 1423 -5 1487 -4
rect 1432 -7 1487 -5
rect 1492 -54 1499 50
rect 1455 -61 1499 -54
rect 1225 -118 1273 -113
rect 1301 -118 1304 -113
rect 1036 -167 1216 -161
rect 1028 -168 1216 -167
rect 1034 -187 1038 -168
rect 1063 -187 1067 -168
rect 1092 -187 1096 -168
rect 1121 -187 1125 -168
rect 1142 -182 1183 -178
rect 1142 -187 1146 -182
rect 1150 -187 1154 -182
rect 1179 -187 1183 -182
rect 1035 -230 1038 -225
rect 1055 -259 1059 -191
rect 1084 -242 1088 -191
rect 1113 -198 1117 -191
rect 1142 -198 1146 -191
rect 1113 -201 1146 -198
rect 1171 -198 1175 -191
rect 1200 -198 1204 -191
rect 1171 -201 1204 -198
rect 1149 -220 1157 -216
rect 1154 -221 1157 -220
rect 1200 -224 1204 -201
rect 1200 -234 1208 -224
rect 1084 -247 1186 -242
rect 1084 -259 1088 -247
rect 1182 -248 1186 -247
rect 1200 -251 1204 -234
rect 1142 -259 1146 -258
rect 1200 -259 1204 -256
rect 1117 -263 1121 -259
rect 1175 -263 1179 -259
rect 1034 -267 1038 -263
rect 1063 -267 1067 -263
rect 1092 -267 1096 -263
rect 1150 -267 1154 -263
rect 996 -274 1219 -267
rect 996 -332 1008 -274
rect 1225 -295 1232 -118
rect 1317 -128 1322 -105
rect 1350 -107 1415 -102
rect 1350 -128 1355 -107
rect 1291 -133 1298 -128
rect 1267 -137 1272 -133
rect 1331 -137 1336 -133
rect 1069 -302 1232 -295
rect 1261 -144 1368 -137
rect 1261 -332 1275 -144
rect 996 -334 1275 -332
rect 1590 -334 1608 182
rect 996 -336 1608 -334
rect 393 -339 1608 -336
rect -833 -340 1608 -339
rect -833 -341 -554 -340
rect -207 -341 1608 -340
rect -207 -344 672 -341
rect 1249 -342 1608 -341
<< m2contact >>
rect -840 224 -833 229
rect -809 234 -803 239
rect -724 234 -719 239
rect -662 220 -653 229
rect -620 224 -613 229
rect -726 196 -721 201
rect -669 198 -664 203
rect -591 234 -585 239
rect -506 234 -501 239
rect -446 220 -437 231
rect -389 226 -382 231
rect -508 196 -503 201
rect -451 198 -446 203
rect -358 236 -352 241
rect -273 236 -268 241
rect -181 222 -172 232
rect -129 227 -122 232
rect -275 198 -270 203
rect -218 200 -213 205
rect -98 237 -92 242
rect -13 237 -8 242
rect 92 224 104 232
rect -15 199 -10 204
rect 42 201 47 206
rect -808 26 -803 31
rect -764 36 -758 41
rect -777 25 -772 30
rect -695 36 -690 41
rect -697 -2 -692 3
rect -640 0 -635 5
rect -868 -168 -854 -154
rect -627 -18 -618 -10
rect -578 21 -573 26
rect -547 21 -542 26
rect -490 32 -482 37
rect -387 15 -382 20
rect -352 19 -344 26
rect -586 -7 -577 1
rect -483 -6 -474 2
rect -440 -61 -430 -54
rect -406 -13 -397 -5
rect -383 -61 -374 -54
rect -534 -118 -528 -112
rect -801 -167 -793 -160
rect -802 -231 -794 -224
rect -770 -220 -764 -215
rect -767 -231 -762 -226
rect -685 -220 -680 -215
rect -687 -258 -682 -253
rect -630 -256 -625 -251
rect -765 -302 -760 -295
rect -182 23 -177 28
rect -138 33 -132 38
rect -151 22 -146 27
rect -69 33 -64 38
rect -71 -5 -66 0
rect -14 -3 -9 2
rect -242 -171 -228 -157
rect -1 -21 8 -13
rect 48 18 53 23
rect 79 18 84 23
rect 136 29 144 34
rect 239 12 244 17
rect 278 16 284 21
rect 40 -10 49 -2
rect 143 -9 152 -1
rect 186 -64 196 -57
rect 220 -16 229 -8
rect 243 -64 252 -57
rect 92 -121 98 -115
rect -175 -170 -167 -163
rect -175 -236 -168 -227
rect -144 -223 -138 -218
rect -141 -234 -136 -229
rect -59 -223 -54 -218
rect -61 -261 -56 -256
rect -4 -259 1 -254
rect -139 -305 -134 -298
rect 418 23 423 28
rect 462 33 468 38
rect 449 22 454 27
rect 531 33 536 38
rect 529 -5 534 0
rect 586 -3 591 2
rect 358 -171 372 -157
rect 599 -21 608 -13
rect 648 18 653 23
rect 679 18 684 23
rect 736 29 744 34
rect 839 12 844 17
rect 878 16 883 21
rect 640 -10 649 -2
rect 743 -9 752 -1
rect 786 -64 796 -57
rect 820 -16 829 -8
rect 843 -64 852 -57
rect 692 -121 698 -115
rect 425 -170 433 -163
rect 425 -233 433 -226
rect 456 -223 462 -218
rect 459 -234 464 -229
rect 541 -223 546 -218
rect 539 -261 544 -256
rect 596 -259 601 -254
rect 461 -305 466 -298
rect 1021 26 1026 31
rect 1065 36 1071 41
rect 1052 25 1057 30
rect 1134 36 1139 41
rect 1132 -2 1137 3
rect 1189 0 1194 5
rect 961 -168 975 -154
rect 1202 -18 1211 -10
rect 1251 21 1256 26
rect 1282 21 1287 26
rect 1339 32 1347 37
rect 1442 15 1447 20
rect 1243 -7 1252 1
rect 1346 -6 1355 2
rect 1389 -61 1399 -54
rect 1423 -13 1432 -5
rect 1446 -61 1455 -54
rect 1295 -118 1301 -112
rect 1028 -167 1036 -160
rect 1028 -231 1035 -224
rect 1059 -220 1065 -215
rect 1062 -231 1067 -226
rect 1144 -220 1149 -215
rect 1142 -258 1147 -253
rect 1199 -256 1204 -251
rect 1064 -302 1069 -295
<< metal2 >>
rect -859 298 -41 304
rect -859 242 -853 298
rect -906 237 -853 242
rect -906 -225 -900 237
rect -859 229 -853 237
rect -803 234 -724 238
rect -620 229 -616 298
rect -585 234 -506 238
rect -389 231 -385 298
rect -352 236 -273 240
rect -129 232 -125 298
rect -92 237 -13 241
rect -859 224 -840 229
rect -437 220 -423 231
rect -721 198 -669 201
rect -658 100 -653 220
rect -503 198 -451 201
rect -427 134 -423 220
rect 104 224 1127 231
rect -270 200 -218 203
rect -181 158 -172 222
rect -10 201 42 204
rect -181 148 457 158
rect -427 131 -95 134
rect -777 97 -543 100
rect -99 97 -95 131
rect 452 97 457 148
rect 1115 100 1122 224
rect 1052 97 1286 100
rect -808 21 -803 26
rect -777 30 -773 97
rect -758 36 -695 40
rect -547 26 -543 97
rect -151 94 83 97
rect -453 61 -382 65
rect -453 37 -449 61
rect -482 32 -449 37
rect -659 21 -578 25
rect -808 18 -655 21
rect -387 20 -382 61
rect -344 19 -298 26
rect -692 0 -640 3
rect -586 -12 -577 -7
rect -618 -18 -577 -12
rect -627 -19 -577 -18
rect -482 -17 -475 -6
rect -406 -17 -397 -13
rect -482 -22 -397 -17
rect -430 -61 -383 -54
rect -854 -167 -801 -162
rect -854 -168 -795 -167
rect -764 -220 -685 -216
rect -906 -231 -802 -225
rect -800 -314 -794 -231
rect -765 -295 -762 -231
rect -682 -256 -630 -253
rect -534 -314 -528 -118
rect -302 -227 -298 19
rect -182 18 -177 23
rect -151 27 -147 94
rect -132 33 -69 37
rect 79 23 83 94
rect 449 94 683 97
rect 173 58 244 62
rect 173 34 177 58
rect 144 29 177 34
rect -33 18 48 22
rect -182 15 -29 18
rect 239 17 244 58
rect 278 21 320 22
rect 284 16 320 21
rect -66 -3 -14 0
rect 40 -15 49 -10
rect 8 -21 49 -15
rect -1 -22 49 -21
rect 144 -20 151 -9
rect 220 -20 229 -16
rect 144 -25 229 -20
rect 196 -64 243 -57
rect -228 -170 -175 -165
rect -228 -171 -169 -170
rect -138 -223 -59 -219
rect -302 -235 -175 -227
rect -800 -318 -528 -314
rect -174 -317 -168 -236
rect -139 -298 -136 -234
rect -56 -259 -4 -256
rect 92 -317 98 -121
rect 316 -227 320 16
rect 418 18 423 23
rect 449 27 453 94
rect 468 33 531 37
rect 679 23 683 94
rect 773 58 844 62
rect 773 34 777 58
rect 744 29 777 34
rect 567 18 648 22
rect 418 15 571 18
rect 839 17 844 58
rect 1021 21 1026 26
rect 1052 30 1056 97
rect 1071 36 1134 40
rect 1282 26 1286 97
rect 1376 61 1447 65
rect 1376 37 1380 61
rect 1347 32 1380 37
rect 1170 21 1251 25
rect 883 16 924 20
rect 1021 18 1174 21
rect 1442 20 1447 61
rect 534 -3 586 0
rect 640 -15 649 -10
rect 608 -21 649 -15
rect 599 -22 649 -21
rect 744 -20 751 -9
rect 820 -20 829 -16
rect 744 -25 829 -20
rect 796 -64 843 -57
rect 372 -170 425 -165
rect 372 -171 431 -170
rect 462 -223 541 -219
rect 316 -233 425 -227
rect -174 -321 98 -317
rect 426 -317 432 -233
rect 461 -298 464 -234
rect 544 -259 596 -256
rect 692 -317 698 -121
rect 914 -224 923 16
rect 1137 0 1189 3
rect 1243 -12 1252 -7
rect 1211 -18 1252 -12
rect 1202 -19 1252 -18
rect 1347 -17 1354 -6
rect 1423 -17 1432 -13
rect 1347 -22 1432 -17
rect 1399 -61 1446 -54
rect 975 -167 1028 -162
rect 975 -168 1034 -167
rect 1065 -220 1144 -216
rect 914 -229 1028 -224
rect 914 -230 923 -229
rect 426 -321 698 -317
rect 1029 -314 1035 -231
rect 1064 -295 1067 -231
rect 1147 -256 1199 -253
rect 1295 -314 1301 -118
rect 1029 -318 1301 -314
<< labels >>
rlabel metal2 -849 226 -849 226 1 node_m
rlabel metal1 -805 224 -805 224 1 node_b0
rlabel metal1 -664 225 -664 225 1 node_z0
rlabel metal1 -584 225 -584 225 1 node_b1
rlabel m2contact -443 224 -443 224 1 node_z1
rlabel metal1 -351 226 -351 226 1 node_b2
rlabel metal1 -94 228 -94 228 1 node_b3
rlabel metal1 -734 288 -734 288 1 vdd
rlabel metal1 -780 183 -780 183 1 gnd
rlabel metal1 1479 20 1479 20 1 node_c
rlabel m2contact -807 28 -807 28 1 node_a0
rlabel m2contact -180 25 -180 25 1 node_a1
rlabel m2contact 420 25 420 25 1 node_a2
rlabel m2contact 1024 28 1024 28 1 node_a3
rlabel metal1 -353 21 -353 21 1 node_c0
rlabel metal1 875 17 875 17 1 node_c2
rlabel m2contact 279 18 279 18 1 node_c1
rlabel metal1 -626 -229 -626 -229 1 node_s0
rlabel metal1 0 -232 0 -232 1 node_s1
rlabel metal1 601 -232 601 -232 1 node_s2
rlabel metal1 1203 -229 1203 -229 1 node_s3
<< end >>
