.include TSMC_180nm.txt
.include not.sub

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param wp1 = wn1
.param lp1 = {LAMBDA}


.global gnd

Vdd node_x gnd 'SUPPLY'

V_in node_in gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 50ns)

X1 node_in node_out node_x gnd not 

C1 node_out gnd 100f

.tran 1n 800n

.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(node_in) v(node_out)+2
hardcopy image.ps v(node_in) v(node_out)+2
.end
.endc