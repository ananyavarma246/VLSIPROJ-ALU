magic
tech scmos
timestamp 1700142763
<< nwell >>
rect 20 162 33 167
rect -251 160 -238 161
rect -308 130 -208 160
rect -172 131 -72 161
rect -37 132 63 162
rect 157 160 170 165
rect 100 130 200 160
rect -252 40 -239 45
rect -106 41 -93 46
rect 24 44 37 49
rect -309 10 -209 40
rect -163 11 -63 41
rect -33 14 67 44
rect 165 43 178 48
rect 108 13 208 43
<< ntransistor >>
rect -293 84 -289 93
rect -261 84 -257 93
rect -227 84 -223 93
rect -157 85 -153 94
rect -125 85 -121 94
rect -91 85 -87 94
rect -22 86 -18 95
rect 10 86 14 95
rect 44 86 48 95
rect 115 84 119 93
rect 147 84 151 93
rect 181 84 185 93
rect -294 -36 -290 -27
rect -262 -36 -258 -27
rect -228 -36 -224 -27
rect -148 -35 -144 -26
rect -116 -35 -112 -26
rect -82 -35 -78 -26
rect -18 -32 -14 -23
rect 14 -32 18 -23
rect 48 -32 52 -23
rect 123 -33 127 -24
rect 155 -33 159 -24
rect 189 -33 193 -24
<< ptransistor >>
rect -293 142 -289 151
rect -261 142 -257 151
rect -227 142 -223 151
rect -157 143 -153 152
rect -125 143 -121 152
rect -91 143 -87 152
rect -22 144 -18 153
rect 10 144 14 153
rect 44 144 48 153
rect 115 142 119 151
rect 147 142 151 151
rect 181 142 185 151
rect -294 22 -290 31
rect -262 22 -258 31
rect -228 22 -224 31
rect -148 23 -144 32
rect -116 23 -112 32
rect -82 23 -78 32
rect -18 26 -14 35
rect 14 26 18 35
rect 48 26 52 35
rect 123 25 127 34
rect 155 25 159 34
rect 189 25 193 34
<< ndiffusion >>
rect -297 88 -293 93
rect -302 84 -293 88
rect -289 88 -283 93
rect -289 84 -278 88
rect -266 88 -261 93
rect -271 84 -261 88
rect -257 88 -252 93
rect -257 84 -247 88
rect -233 88 -227 93
rect -238 84 -227 88
rect -223 88 -219 93
rect -223 84 -214 88
rect -161 89 -157 94
rect -166 85 -157 89
rect -153 89 -147 94
rect -153 85 -142 89
rect -130 89 -125 94
rect -135 85 -125 89
rect -121 89 -116 94
rect -121 85 -111 89
rect -97 89 -91 94
rect -102 85 -91 89
rect -87 89 -83 94
rect -87 85 -78 89
rect -26 90 -22 95
rect -31 86 -22 90
rect -18 90 -12 95
rect -18 86 -7 90
rect 5 90 10 95
rect 0 86 10 90
rect 14 90 19 95
rect 14 86 24 90
rect 38 90 44 95
rect 33 86 44 90
rect 48 90 52 95
rect 48 86 57 90
rect 111 88 115 93
rect 106 84 115 88
rect 119 88 125 93
rect 119 84 130 88
rect 142 88 147 93
rect 137 84 147 88
rect 151 88 156 93
rect 151 84 161 88
rect 175 88 181 93
rect 170 84 181 88
rect 185 88 189 93
rect 185 84 194 88
rect -298 -32 -294 -27
rect -303 -36 -294 -32
rect -290 -32 -284 -27
rect -290 -36 -279 -32
rect -267 -32 -262 -27
rect -272 -36 -262 -32
rect -258 -32 -253 -27
rect -258 -36 -248 -32
rect -234 -32 -228 -27
rect -239 -36 -228 -32
rect -224 -32 -220 -27
rect -224 -36 -215 -32
rect -152 -31 -148 -26
rect -157 -35 -148 -31
rect -144 -31 -138 -26
rect -144 -35 -133 -31
rect -121 -31 -116 -26
rect -126 -35 -116 -31
rect -112 -31 -107 -26
rect -112 -35 -102 -31
rect -88 -31 -82 -26
rect -93 -35 -82 -31
rect -78 -31 -74 -26
rect -78 -35 -69 -31
rect -22 -28 -18 -23
rect -27 -32 -18 -28
rect -14 -28 -8 -23
rect -14 -32 -3 -28
rect 9 -28 14 -23
rect 4 -32 14 -28
rect 18 -28 23 -23
rect 18 -32 28 -28
rect 42 -28 48 -23
rect 37 -32 48 -28
rect 52 -28 56 -23
rect 52 -32 61 -28
rect 119 -29 123 -24
rect 114 -33 123 -29
rect 127 -29 133 -24
rect 127 -33 138 -29
rect 150 -29 155 -24
rect 145 -33 155 -29
rect 159 -29 164 -24
rect 159 -33 169 -29
rect 183 -29 189 -24
rect 178 -33 189 -29
rect 193 -29 197 -24
rect 193 -33 202 -29
<< pdiffusion >>
rect -297 146 -293 151
rect -302 142 -293 146
rect -289 146 -283 151
rect -289 142 -278 146
rect -266 146 -261 151
rect -271 142 -261 146
rect -257 146 -252 151
rect -257 142 -247 146
rect -233 146 -227 151
rect -238 142 -227 146
rect -223 146 -219 151
rect -223 142 -214 146
rect -161 147 -157 152
rect -166 143 -157 147
rect -153 147 -147 152
rect -153 143 -142 147
rect -130 147 -125 152
rect -135 143 -125 147
rect -121 147 -116 152
rect -121 143 -111 147
rect -97 147 -91 152
rect -102 143 -91 147
rect -87 147 -83 152
rect -87 143 -78 147
rect -26 148 -22 153
rect -31 144 -22 148
rect -18 148 -12 153
rect -18 144 -7 148
rect 5 148 10 153
rect 0 144 10 148
rect 14 148 19 153
rect 14 144 24 148
rect 38 148 44 153
rect 33 144 44 148
rect 48 148 52 153
rect 48 144 57 148
rect 111 146 115 151
rect 106 142 115 146
rect 119 146 125 151
rect 119 142 130 146
rect 142 146 147 151
rect 137 142 147 146
rect 151 146 156 151
rect 151 142 161 146
rect 175 146 181 151
rect 170 142 181 146
rect 185 146 189 151
rect 185 142 194 146
rect -298 26 -294 31
rect -303 22 -294 26
rect -290 26 -284 31
rect -290 22 -279 26
rect -267 26 -262 31
rect -272 22 -262 26
rect -258 26 -253 31
rect -258 22 -248 26
rect -234 26 -228 31
rect -239 22 -228 26
rect -224 26 -220 31
rect -224 22 -215 26
rect -152 27 -148 32
rect -157 23 -148 27
rect -144 27 -138 32
rect -144 23 -133 27
rect -121 27 -116 32
rect -126 23 -116 27
rect -112 27 -107 32
rect -112 23 -102 27
rect -88 27 -82 32
rect -93 23 -82 27
rect -78 27 -74 32
rect -78 23 -69 27
rect -22 30 -18 35
rect -27 26 -18 30
rect -14 30 -8 35
rect -14 26 -3 30
rect 9 30 14 35
rect 4 26 14 30
rect 18 30 23 35
rect 18 26 28 30
rect 42 30 48 35
rect 37 26 48 30
rect 52 30 56 35
rect 52 26 61 30
rect 119 29 123 34
rect 114 25 123 29
rect 127 29 133 34
rect 127 25 138 29
rect 150 29 155 34
rect 145 25 155 29
rect 159 29 164 34
rect 159 25 169 29
rect 183 29 189 34
rect 178 25 189 29
rect 193 29 197 34
rect 193 25 202 29
<< ndcontact >>
rect -302 88 -297 93
rect -283 88 -278 93
rect -271 88 -266 93
rect -252 88 -247 93
rect -238 88 -233 93
rect -219 88 -214 93
rect -166 89 -161 94
rect -147 89 -142 94
rect -135 89 -130 94
rect -116 89 -111 94
rect -102 89 -97 94
rect -83 89 -78 94
rect -31 90 -26 95
rect -12 90 -7 95
rect 0 90 5 95
rect 19 90 24 95
rect 33 90 38 95
rect 52 90 57 95
rect 106 88 111 93
rect 125 88 130 93
rect 137 88 142 93
rect 156 88 161 93
rect 170 88 175 93
rect 189 88 194 93
rect -303 -32 -298 -27
rect -284 -32 -279 -27
rect -272 -32 -267 -27
rect -253 -32 -248 -27
rect -239 -32 -234 -27
rect -220 -32 -215 -27
rect -157 -31 -152 -26
rect -138 -31 -133 -26
rect -126 -31 -121 -26
rect -107 -31 -102 -26
rect -93 -31 -88 -26
rect -74 -31 -69 -26
rect -27 -28 -22 -23
rect -8 -28 -3 -23
rect 4 -28 9 -23
rect 23 -28 28 -23
rect 37 -28 42 -23
rect 56 -28 61 -23
rect 114 -29 119 -24
rect 133 -29 138 -24
rect 145 -29 150 -24
rect 164 -29 169 -24
rect 178 -29 183 -24
rect 197 -29 202 -24
<< pdcontact >>
rect -302 146 -297 151
rect -283 146 -278 151
rect -271 146 -266 151
rect -252 146 -247 151
rect -238 146 -233 151
rect -219 146 -214 151
rect -166 147 -161 152
rect -147 147 -142 152
rect -135 147 -130 152
rect -116 147 -111 152
rect -102 147 -97 152
rect -83 147 -78 152
rect -31 148 -26 153
rect -12 148 -7 153
rect 0 148 5 153
rect 19 148 24 153
rect 33 148 38 153
rect 52 148 57 153
rect 106 146 111 151
rect 125 146 130 151
rect 137 146 142 151
rect 156 146 161 151
rect 170 146 175 151
rect 189 146 194 151
rect -303 26 -298 31
rect -284 26 -279 31
rect -272 26 -267 31
rect -253 26 -248 31
rect -239 26 -234 31
rect -220 26 -215 31
rect -157 27 -152 32
rect -138 27 -133 32
rect -126 27 -121 32
rect -107 27 -102 32
rect -93 27 -88 32
rect -74 27 -69 32
rect -27 30 -22 35
rect -8 30 -3 35
rect 4 30 9 35
rect 23 30 28 35
rect 37 30 42 35
rect 56 30 61 35
rect 114 29 119 34
rect 133 29 138 34
rect 145 29 150 34
rect 164 29 169 34
rect 178 29 183 34
rect 197 29 202 34
<< polysilicon >>
rect -293 151 -289 157
rect -261 151 -257 155
rect -227 151 -223 155
rect -157 152 -153 158
rect -125 152 -121 156
rect -91 152 -87 156
rect -22 153 -18 159
rect 10 153 14 157
rect 44 153 48 157
rect 115 151 119 157
rect 147 151 151 155
rect 181 151 185 155
rect -293 108 -289 142
rect -292 103 -289 108
rect -293 93 -289 103
rect -261 93 -257 142
rect -227 93 -223 142
rect -157 109 -153 143
rect -156 104 -153 109
rect -157 94 -153 104
rect -125 94 -121 143
rect -91 94 -87 143
rect -22 110 -18 144
rect -21 105 -18 110
rect -22 95 -18 105
rect 10 95 14 144
rect 44 95 48 144
rect 115 108 119 142
rect 116 103 119 108
rect 115 93 119 103
rect 147 93 151 142
rect 181 93 185 142
rect -293 81 -289 84
rect -261 81 -257 84
rect -227 81 -223 84
rect -157 82 -153 85
rect -125 82 -121 85
rect -91 82 -87 85
rect -22 83 -18 86
rect 10 83 14 86
rect 44 83 48 86
rect 115 81 119 84
rect 147 81 151 84
rect 181 81 185 84
rect -294 31 -290 37
rect -262 31 -258 35
rect -228 31 -224 35
rect -148 32 -144 38
rect -116 32 -112 36
rect -82 32 -78 36
rect -18 35 -14 41
rect 14 35 18 39
rect 48 35 52 39
rect 123 34 127 40
rect 155 34 159 38
rect 189 34 193 38
rect -294 -12 -290 22
rect -293 -17 -290 -12
rect -294 -27 -290 -17
rect -262 -27 -258 22
rect -228 -27 -224 22
rect -148 -11 -144 23
rect -147 -16 -144 -11
rect -148 -26 -144 -16
rect -116 -26 -112 23
rect -82 -26 -78 23
rect -18 -8 -14 26
rect -17 -13 -14 -8
rect -18 -23 -14 -13
rect 14 -23 18 26
rect 48 -23 52 26
rect 123 -9 127 25
rect 124 -14 127 -9
rect 123 -24 127 -14
rect 155 -24 159 25
rect 189 -24 193 25
rect -18 -35 -14 -32
rect 14 -35 18 -32
rect 48 -35 52 -32
rect -294 -39 -290 -36
rect -262 -39 -258 -36
rect -228 -39 -224 -36
rect -148 -38 -144 -35
rect -116 -38 -112 -35
rect -82 -38 -78 -35
rect 123 -36 127 -33
rect 155 -36 159 -33
rect 189 -36 193 -33
<< polycontact >>
rect -296 103 -292 108
rect -265 103 -261 108
rect -233 116 -227 122
rect -160 104 -156 109
rect -129 104 -125 109
rect -97 117 -91 123
rect -25 105 -21 110
rect 6 105 10 110
rect 38 118 44 124
rect 112 103 116 108
rect 143 103 147 108
rect 175 116 181 122
rect -297 -17 -293 -12
rect -266 -17 -262 -12
rect -234 -4 -228 2
rect -151 -16 -147 -11
rect -120 -16 -116 -11
rect -88 -3 -82 3
rect -21 -13 -17 -8
rect 10 -13 14 -8
rect 42 0 48 6
rect 120 -14 124 -9
rect 151 -14 155 -9
rect 183 -1 189 5
<< metal1 >>
rect -335 167 -70 168
rect -38 167 65 169
rect -335 162 202 167
rect -335 161 -70 162
rect -449 83 -422 93
rect -334 47 -329 161
rect -309 160 -206 161
rect -302 151 -297 160
rect -271 151 -266 160
rect -238 151 -233 160
rect -166 152 -161 161
rect -135 152 -130 161
rect -102 152 -97 161
rect -31 153 -26 162
rect 0 153 5 162
rect 33 153 38 162
rect 85 161 202 162
rect 99 160 202 161
rect -283 122 -278 146
rect -252 122 -247 146
rect -283 116 -233 122
rect -219 119 -214 146
rect -147 123 -142 147
rect -116 123 -111 147
rect -305 103 -296 108
rect -269 103 -265 108
rect -252 93 -247 116
rect -219 114 -211 119
rect -147 117 -97 123
rect -83 120 -78 147
rect -12 124 -7 148
rect 19 124 24 148
rect -219 93 -214 114
rect -169 104 -160 109
rect -131 104 -129 109
rect -116 94 -111 117
rect -83 115 -75 120
rect -12 118 38 124
rect 52 121 57 148
rect 106 151 111 160
rect 137 151 142 160
rect 170 151 175 160
rect 125 122 130 146
rect 156 122 161 146
rect -83 94 -78 115
rect -34 105 -25 110
rect 4 105 6 110
rect 19 95 24 118
rect 52 116 60 121
rect 125 116 175 122
rect 189 119 194 146
rect 52 95 57 116
rect 103 103 112 108
rect 141 103 143 108
rect -278 88 -271 93
rect -142 89 -135 94
rect -7 90 0 95
rect 156 93 161 116
rect 189 114 197 119
rect 189 93 194 114
rect -302 84 -297 88
rect -238 84 -233 88
rect -166 85 -161 89
rect -102 85 -97 89
rect -31 86 -26 90
rect 33 86 38 90
rect 130 88 137 93
rect -172 84 -59 85
rect -37 84 76 86
rect 106 84 111 88
rect 170 84 175 88
rect -308 83 -195 84
rect -172 83 238 84
rect -308 82 238 83
rect -309 79 238 82
rect -308 78 -52 79
rect -308 77 -195 78
rect 100 77 238 79
rect -34 50 69 51
rect -65 48 210 50
rect -334 45 -207 47
rect -164 45 210 48
rect -334 44 210 45
rect -334 42 -61 44
rect -334 40 -207 42
rect -164 41 -61 42
rect -303 31 -298 40
rect -272 31 -267 40
rect -239 31 -234 40
rect -157 32 -152 41
rect -126 32 -121 41
rect -93 32 -88 41
rect -27 35 -22 44
rect 4 35 9 44
rect 37 35 42 44
rect 107 43 210 44
rect -284 2 -279 26
rect -253 2 -248 26
rect -284 -4 -234 2
rect -220 -1 -215 26
rect -138 3 -133 27
rect -107 3 -102 27
rect -306 -17 -297 -12
rect -268 -17 -266 -12
rect -253 -27 -248 -4
rect -220 -6 -212 -1
rect -138 -3 -88 3
rect -74 0 -69 27
rect -8 6 -3 30
rect 23 6 28 30
rect -8 0 42 6
rect 56 3 61 30
rect 114 34 119 43
rect 145 34 150 43
rect 178 34 183 43
rect 133 5 138 29
rect 164 5 169 29
rect -220 -27 -215 -6
rect -160 -16 -151 -11
rect -123 -16 -120 -11
rect -107 -26 -102 -3
rect -74 -5 -66 0
rect -74 -26 -69 -5
rect -30 -13 -21 -8
rect 6 -13 10 -8
rect 23 -23 28 0
rect 56 -2 64 3
rect 133 -1 183 5
rect 197 2 202 29
rect 56 -23 61 -2
rect 111 -14 120 -9
rect 147 -14 151 -9
rect -279 -32 -272 -27
rect -133 -31 -126 -26
rect -3 -28 4 -23
rect 164 -24 169 -1
rect 197 -3 205 2
rect 197 -24 202 -3
rect -303 -36 -298 -32
rect -239 -36 -234 -32
rect -157 -35 -152 -31
rect -93 -35 -88 -31
rect -27 -32 -22 -28
rect 37 -32 42 -28
rect 138 -29 145 -24
rect -33 -34 80 -32
rect 114 -33 119 -29
rect 178 -33 183 -29
rect 230 -33 238 77
rect -63 -35 80 -34
rect 108 -35 238 -33
rect -202 -36 238 -35
rect -324 -38 238 -36
rect -324 -39 80 -38
rect -324 -42 -29 -39
rect 108 -40 238 -38
rect -324 -43 -162 -42
<< m2contact >>
rect -422 83 -408 93
rect -274 103 -269 108
rect -136 104 -131 109
rect -1 105 4 110
rect 136 103 141 108
rect -273 -17 -268 -12
rect -128 -16 -123 -11
rect 1 -13 6 -8
rect 142 -14 147 -9
<< metal2 >>
rect -405 181 239 192
rect -405 93 -395 181
rect -274 108 -269 181
rect -136 109 -131 181
rect -1 110 4 181
rect 136 108 141 181
rect -408 83 -395 93
rect -406 -55 -395 83
rect -273 -55 -268 -17
rect -128 -55 -123 -16
rect 1 -55 6 -13
rect 142 -55 147 -14
rect -406 -63 267 -55
<< labels >>
rlabel metal1 -174 164 -174 164 5 vdd
rlabel metal1 -175 -40 -175 -40 1 gnd
rlabel metal1 -302 -16 -302 -16 1 node_bo
rlabel metal1 -153 -13 -153 -13 1 node_b1
rlabel metal1 -26 -11 -26 -11 1 node_b2
rlabel metal1 116 -12 116 -12 1 node_b3
rlabel metal1 -300 106 -300 106 1 node_a0
rlabel metal1 -164 106 -164 106 1 node_a1
rlabel metal1 -29 107 -29 107 1 node_a2
rlabel metal1 106 104 106 104 1 node_a3
rlabel metal1 -214 116 -214 116 1 node_c0
rlabel metal1 -77 116 -77 116 1 node_c1
rlabel metal1 59 118 59 118 1 node_c2
rlabel metal1 196 117 196 117 1 node_c3
rlabel metal1 -214 -3 -214 -3 1 node_d0
rlabel metal1 -68 -3 -68 -3 1 node_d1
rlabel metal1 63 -1 63 -1 1 node_d2
rlabel metal1 202 0 202 0 1 node_d3
rlabel metal1 -440 87 -440 87 1 enable
<< end >>
