magic
tech scmos
timestamp 1699688820
<< nwell >>
rect -117 206 -47 222
<< ntransistor >>
rect -102 171 -100 175
rect -84 171 -82 175
rect -65 171 -63 175
<< ptransistor >>
rect -102 212 -100 216
rect -84 212 -82 216
rect -65 212 -63 216
<< ndiffusion >>
rect -104 171 -102 175
rect -100 171 -98 175
rect -86 171 -84 175
rect -82 171 -80 175
rect -67 171 -65 175
rect -63 171 -61 175
<< pdiffusion >>
rect -104 212 -102 216
rect -100 212 -98 216
rect -86 212 -84 216
rect -82 212 -80 216
rect -67 212 -65 216
rect -63 212 -61 216
<< ndcontact >>
rect -108 171 -104 175
rect -98 171 -94 175
rect -90 171 -86 175
rect -80 171 -76 175
rect -71 171 -67 175
rect -61 171 -57 175
<< pdcontact >>
rect -108 212 -104 216
rect -98 212 -94 216
rect -90 212 -86 216
rect -80 212 -76 216
rect -71 212 -67 216
rect -61 212 -57 216
<< polysilicon >>
rect -102 216 -100 219
rect -84 216 -82 219
rect -65 216 -63 219
rect -102 189 -100 212
rect -84 191 -82 212
rect -65 192 -63 212
rect -101 185 -100 189
rect -83 187 -82 191
rect -64 188 -63 192
rect -102 175 -100 185
rect -84 175 -82 187
rect -65 175 -63 188
rect -102 168 -100 171
rect -84 168 -82 171
rect -65 168 -63 171
<< polycontact >>
rect -105 185 -101 189
rect -87 187 -83 191
rect -68 188 -64 192
<< metal1 >>
rect -122 222 -46 227
rect -108 216 -104 222
rect -71 216 -67 222
rect -94 212 -90 216
rect -80 192 -76 212
rect -61 195 -57 212
rect -108 185 -105 189
rect -89 187 -87 191
rect -80 188 -68 192
rect -61 191 -52 195
rect -80 183 -76 188
rect -98 180 -76 183
rect -98 175 -94 180
rect -80 175 -76 180
rect -61 175 -57 191
rect -108 168 -104 171
rect -90 168 -86 171
rect -71 168 -67 171
rect -112 165 -48 168
<< labels >>
rlabel metal1 -90 225 -90 225 5 vdd
rlabel metal1 -107 187 -107 187 1 node_a
rlabel metal1 -88 190 -88 190 1 node_b
rlabel metal1 -71 191 -71 191 1 node_inter
rlabel metal1 -56 194 -56 194 1 node_out
rlabel metal1 -88 166 -88 166 1 gnd
rlabel metal1 -93 214 -93 214 1 node_x
<< end >>
