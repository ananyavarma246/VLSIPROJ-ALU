magic
tech scmos
timestamp 1700167176
<< nwell >>
rect -1105 547 -901 579
rect -1106 300 -902 332
rect -752 244 -477 285
rect -1102 74 -898 106
rect -1105 -133 -901 -101
<< ntransistor >>
rect -1089 472 -1086 478
rect -1054 472 -1051 478
rect -1019 472 -1016 478
rect -987 472 -984 478
rect -956 472 -953 478
rect -923 472 -920 478
rect -1090 225 -1087 231
rect -1055 225 -1052 231
rect -1020 225 -1017 231
rect -988 225 -985 231
rect -957 225 -954 231
rect -924 225 -921 231
rect -730 160 -726 171
rect -684 160 -680 171
rect -639 160 -635 171
rect -596 160 -592 171
rect -551 160 -547 171
rect -508 160 -504 171
rect -1086 -1 -1083 5
rect -1051 -1 -1048 5
rect -1016 -1 -1013 5
rect -984 -1 -981 5
rect -953 -1 -950 5
rect -920 -1 -917 5
rect -1089 -208 -1086 -202
rect -1054 -208 -1051 -202
rect -1019 -208 -1016 -202
rect -987 -208 -984 -202
rect -956 -208 -953 -202
rect -923 -208 -920 -202
<< ptransistor >>
rect -1089 561 -1086 567
rect -1054 561 -1051 567
rect -1019 561 -1016 567
rect -987 561 -984 567
rect -956 561 -953 567
rect -923 561 -920 567
rect -1090 314 -1087 320
rect -1055 314 -1052 320
rect -1020 314 -1017 320
rect -988 314 -985 320
rect -957 314 -954 320
rect -924 314 -921 320
rect -730 263 -726 274
rect -684 263 -680 274
rect -639 263 -635 274
rect -596 263 -592 274
rect -551 263 -547 274
rect -508 263 -504 274
rect -1086 88 -1083 94
rect -1051 88 -1048 94
rect -1016 88 -1013 94
rect -984 88 -981 94
rect -953 88 -950 94
rect -920 88 -917 94
rect -1089 -119 -1086 -113
rect -1054 -119 -1051 -113
rect -1019 -119 -1016 -113
rect -987 -119 -984 -113
rect -956 -119 -953 -113
rect -923 -119 -920 -113
<< ndiffusion >>
rect -1095 474 -1089 478
rect -1099 472 -1089 474
rect -1086 474 -1076 478
rect -1086 472 -1072 474
rect -1061 474 -1054 478
rect -1065 472 -1054 474
rect -1051 474 -1042 478
rect -1051 472 -1038 474
rect -1028 474 -1019 478
rect -1032 472 -1019 474
rect -1016 474 -1009 478
rect -1016 472 -1005 474
rect -996 474 -987 478
rect -1000 472 -987 474
rect -984 474 -977 478
rect -984 472 -973 474
rect -964 474 -956 478
rect -968 472 -956 474
rect -953 474 -945 478
rect -953 472 -941 474
rect -932 474 -923 478
rect -936 472 -923 474
rect -920 474 -913 478
rect -920 472 -909 474
rect -1096 227 -1090 231
rect -1100 225 -1090 227
rect -1087 227 -1077 231
rect -1087 225 -1073 227
rect -1062 227 -1055 231
rect -1066 225 -1055 227
rect -1052 227 -1043 231
rect -1052 225 -1039 227
rect -1029 227 -1020 231
rect -1033 225 -1020 227
rect -1017 227 -1010 231
rect -1017 225 -1006 227
rect -997 227 -988 231
rect -1001 225 -988 227
rect -985 227 -978 231
rect -985 225 -974 227
rect -965 227 -957 231
rect -969 225 -957 227
rect -954 227 -946 231
rect -954 225 -942 227
rect -933 227 -924 231
rect -937 225 -924 227
rect -921 227 -914 231
rect -921 225 -910 227
rect -742 167 -730 171
rect -746 160 -730 167
rect -726 167 -710 171
rect -726 160 -706 167
rect -698 167 -684 171
rect -702 160 -684 167
rect -680 167 -666 171
rect -680 160 -662 167
rect -654 167 -639 171
rect -658 160 -639 167
rect -635 167 -622 171
rect -635 160 -618 167
rect -610 167 -596 171
rect -614 160 -596 167
rect -592 167 -578 171
rect -592 160 -574 167
rect -566 167 -551 171
rect -570 160 -551 167
rect -547 167 -534 171
rect -547 160 -530 167
rect -522 167 -508 171
rect -526 160 -508 167
rect -504 167 -490 171
rect -504 160 -486 167
rect -1092 1 -1086 5
rect -1096 -1 -1086 1
rect -1083 1 -1073 5
rect -1083 -1 -1069 1
rect -1058 1 -1051 5
rect -1062 -1 -1051 1
rect -1048 1 -1039 5
rect -1048 -1 -1035 1
rect -1025 1 -1016 5
rect -1029 -1 -1016 1
rect -1013 1 -1006 5
rect -1013 -1 -1002 1
rect -993 1 -984 5
rect -997 -1 -984 1
rect -981 1 -974 5
rect -981 -1 -970 1
rect -961 1 -953 5
rect -965 -1 -953 1
rect -950 1 -942 5
rect -950 -1 -938 1
rect -929 1 -920 5
rect -933 -1 -920 1
rect -917 1 -910 5
rect -917 -1 -906 1
rect -1095 -206 -1089 -202
rect -1099 -208 -1089 -206
rect -1086 -206 -1076 -202
rect -1086 -208 -1072 -206
rect -1061 -206 -1054 -202
rect -1065 -208 -1054 -206
rect -1051 -206 -1042 -202
rect -1051 -208 -1038 -206
rect -1028 -206 -1019 -202
rect -1032 -208 -1019 -206
rect -1016 -206 -1009 -202
rect -1016 -208 -1005 -206
rect -996 -206 -987 -202
rect -1000 -208 -987 -206
rect -984 -206 -977 -202
rect -984 -208 -973 -206
rect -964 -206 -956 -202
rect -968 -208 -956 -206
rect -953 -206 -945 -202
rect -953 -208 -941 -206
rect -932 -206 -923 -202
rect -936 -208 -923 -206
rect -920 -206 -913 -202
rect -920 -208 -909 -206
<< pdiffusion >>
rect -1095 563 -1089 567
rect -1099 561 -1089 563
rect -1086 563 -1076 567
rect -1086 561 -1072 563
rect -1061 563 -1054 567
rect -1065 561 -1054 563
rect -1051 563 -1042 567
rect -1051 561 -1038 563
rect -1028 563 -1019 567
rect -1032 561 -1019 563
rect -1016 563 -1009 567
rect -1016 561 -1005 563
rect -996 563 -987 567
rect -1000 561 -987 563
rect -984 563 -977 567
rect -984 561 -973 563
rect -964 563 -956 567
rect -968 561 -956 563
rect -953 563 -945 567
rect -953 561 -941 563
rect -932 563 -923 567
rect -936 561 -923 563
rect -920 563 -913 567
rect -920 561 -909 563
rect -1096 316 -1090 320
rect -1100 314 -1090 316
rect -1087 316 -1077 320
rect -1087 314 -1073 316
rect -1062 316 -1055 320
rect -1066 314 -1055 316
rect -1052 316 -1043 320
rect -1052 314 -1039 316
rect -1029 316 -1020 320
rect -1033 314 -1020 316
rect -1017 316 -1010 320
rect -1017 314 -1006 316
rect -997 316 -988 320
rect -1001 314 -988 316
rect -985 316 -978 320
rect -985 314 -974 316
rect -965 316 -957 320
rect -969 314 -957 316
rect -954 316 -946 320
rect -954 314 -942 316
rect -933 316 -924 320
rect -937 314 -924 316
rect -921 316 -914 320
rect -921 314 -910 316
rect -742 270 -730 274
rect -746 263 -730 270
rect -726 270 -710 274
rect -726 263 -706 270
rect -698 270 -684 274
rect -702 263 -684 270
rect -680 270 -666 274
rect -680 263 -662 270
rect -654 270 -639 274
rect -658 263 -639 270
rect -635 270 -622 274
rect -635 263 -618 270
rect -610 270 -596 274
rect -614 263 -596 270
rect -592 270 -578 274
rect -592 263 -574 270
rect -566 270 -551 274
rect -570 263 -551 270
rect -547 270 -534 274
rect -547 263 -530 270
rect -522 270 -508 274
rect -526 263 -508 270
rect -504 270 -490 274
rect -504 263 -486 270
rect -1092 90 -1086 94
rect -1096 88 -1086 90
rect -1083 90 -1073 94
rect -1083 88 -1069 90
rect -1058 90 -1051 94
rect -1062 88 -1051 90
rect -1048 90 -1039 94
rect -1048 88 -1035 90
rect -1025 90 -1016 94
rect -1029 88 -1016 90
rect -1013 90 -1006 94
rect -1013 88 -1002 90
rect -993 90 -984 94
rect -997 88 -984 90
rect -981 90 -974 94
rect -981 88 -970 90
rect -961 90 -953 94
rect -965 88 -953 90
rect -950 90 -942 94
rect -950 88 -938 90
rect -929 90 -920 94
rect -933 88 -920 90
rect -917 90 -910 94
rect -917 88 -906 90
rect -1095 -117 -1089 -113
rect -1099 -119 -1089 -117
rect -1086 -117 -1076 -113
rect -1086 -119 -1072 -117
rect -1061 -117 -1054 -113
rect -1065 -119 -1054 -117
rect -1051 -117 -1042 -113
rect -1051 -119 -1038 -117
rect -1028 -117 -1019 -113
rect -1032 -119 -1019 -117
rect -1016 -117 -1009 -113
rect -1016 -119 -1005 -117
rect -996 -117 -987 -113
rect -1000 -119 -987 -117
rect -984 -117 -977 -113
rect -984 -119 -973 -117
rect -964 -117 -956 -113
rect -968 -119 -956 -117
rect -953 -117 -945 -113
rect -953 -119 -941 -117
rect -932 -117 -923 -113
rect -936 -119 -923 -117
rect -920 -117 -913 -113
rect -920 -119 -909 -117
<< ndcontact >>
rect -1099 474 -1095 478
rect -1076 474 -1072 478
rect -1065 474 -1061 478
rect -1042 474 -1038 478
rect -1032 474 -1028 478
rect -1009 474 -1005 478
rect -1000 474 -996 478
rect -977 474 -973 478
rect -968 474 -964 478
rect -945 474 -941 478
rect -936 474 -932 478
rect -913 474 -909 478
rect -1100 227 -1096 231
rect -1077 227 -1073 231
rect -1066 227 -1062 231
rect -1043 227 -1039 231
rect -1033 227 -1029 231
rect -1010 227 -1006 231
rect -1001 227 -997 231
rect -978 227 -974 231
rect -969 227 -965 231
rect -946 227 -942 231
rect -937 227 -933 231
rect -914 227 -910 231
rect -746 167 -742 171
rect -710 167 -706 171
rect -702 167 -698 171
rect -666 167 -662 171
rect -658 167 -654 171
rect -622 167 -618 171
rect -614 167 -610 171
rect -578 167 -574 171
rect -570 167 -566 171
rect -534 167 -530 171
rect -526 167 -522 171
rect -490 167 -486 171
rect -1096 1 -1092 5
rect -1073 1 -1069 5
rect -1062 1 -1058 5
rect -1039 1 -1035 5
rect -1029 1 -1025 5
rect -1006 1 -1002 5
rect -997 1 -993 5
rect -974 1 -970 5
rect -965 1 -961 5
rect -942 1 -938 5
rect -933 1 -929 5
rect -910 1 -906 5
rect -1099 -206 -1095 -202
rect -1076 -206 -1072 -202
rect -1065 -206 -1061 -202
rect -1042 -206 -1038 -202
rect -1032 -206 -1028 -202
rect -1009 -206 -1005 -202
rect -1000 -206 -996 -202
rect -977 -206 -973 -202
rect -968 -206 -964 -202
rect -945 -206 -941 -202
rect -936 -206 -932 -202
rect -913 -206 -909 -202
<< pdcontact >>
rect -1099 563 -1095 567
rect -1076 563 -1072 567
rect -1065 563 -1061 567
rect -1042 563 -1038 567
rect -1032 563 -1028 567
rect -1009 563 -1005 567
rect -1000 563 -996 567
rect -977 563 -973 567
rect -968 563 -964 567
rect -945 563 -941 567
rect -936 563 -932 567
rect -913 563 -909 567
rect -1100 316 -1096 320
rect -1077 316 -1073 320
rect -1066 316 -1062 320
rect -1043 316 -1039 320
rect -1033 316 -1029 320
rect -1010 316 -1006 320
rect -1001 316 -997 320
rect -978 316 -974 320
rect -969 316 -965 320
rect -946 316 -942 320
rect -937 316 -933 320
rect -914 316 -910 320
rect -746 270 -742 274
rect -710 270 -706 274
rect -702 270 -698 274
rect -666 270 -662 274
rect -658 270 -654 274
rect -622 270 -618 274
rect -614 270 -610 274
rect -578 270 -574 274
rect -570 270 -566 274
rect -534 270 -530 274
rect -526 270 -522 274
rect -490 270 -486 274
rect -1096 90 -1092 94
rect -1073 90 -1069 94
rect -1062 90 -1058 94
rect -1039 90 -1035 94
rect -1029 90 -1025 94
rect -1006 90 -1002 94
rect -997 90 -993 94
rect -974 90 -970 94
rect -965 90 -961 94
rect -942 90 -938 94
rect -933 90 -929 94
rect -910 90 -906 94
rect -1099 -117 -1095 -113
rect -1076 -117 -1072 -113
rect -1065 -117 -1061 -113
rect -1042 -117 -1038 -113
rect -1032 -117 -1028 -113
rect -1009 -117 -1005 -113
rect -1000 -117 -996 -113
rect -977 -117 -973 -113
rect -968 -117 -964 -113
rect -945 -117 -941 -113
rect -936 -117 -932 -113
rect -913 -117 -909 -113
<< polysilicon >>
rect -1054 593 -953 596
rect -1089 567 -1086 576
rect -1054 567 -1051 593
rect -1019 567 -1016 576
rect -987 567 -984 576
rect -956 567 -953 593
rect -923 567 -920 576
rect -1089 478 -1086 561
rect -1054 478 -1051 561
rect -1019 478 -1016 561
rect -987 478 -984 561
rect -956 478 -953 561
rect -923 478 -920 561
rect -1089 461 -1086 472
rect -1054 464 -1051 472
rect -1019 461 -1016 472
rect -987 464 -984 472
rect -956 464 -953 472
rect -923 464 -920 472
rect -1089 459 -1016 461
rect -1055 346 -954 349
rect -1090 320 -1087 329
rect -1055 320 -1052 346
rect -1020 320 -1017 329
rect -988 320 -985 329
rect -957 320 -954 346
rect -924 320 -921 329
rect -1090 231 -1087 314
rect -1055 231 -1052 314
rect -1020 231 -1017 314
rect -988 231 -985 314
rect -957 231 -954 314
rect -924 231 -921 314
rect -730 274 -726 279
rect -684 274 -680 279
rect -639 274 -635 279
rect -596 274 -592 279
rect -551 274 -547 279
rect -508 274 -504 279
rect -1090 214 -1087 225
rect -1055 217 -1052 225
rect -1020 214 -1017 225
rect -988 217 -985 225
rect -957 217 -954 225
rect -924 217 -921 225
rect -1090 212 -1017 214
rect -730 171 -726 263
rect -684 216 -680 263
rect -685 207 -680 216
rect -639 215 -635 263
rect -596 215 -592 263
rect -684 171 -680 207
rect -637 206 -635 215
rect -594 206 -592 215
rect -551 213 -547 263
rect -639 171 -635 206
rect -596 171 -592 206
rect -550 204 -547 213
rect -551 171 -547 204
rect -508 171 -504 263
rect -730 153 -726 160
rect -684 153 -680 160
rect -639 153 -635 160
rect -596 153 -592 160
rect -551 153 -547 160
rect -508 153 -504 160
rect -1051 120 -950 123
rect -1086 94 -1083 103
rect -1051 94 -1048 120
rect -1016 94 -1013 103
rect -984 94 -981 103
rect -953 94 -950 120
rect -920 94 -917 103
rect -1086 5 -1083 88
rect -1051 5 -1048 88
rect -1016 5 -1013 88
rect -984 5 -981 88
rect -953 5 -950 88
rect -920 5 -917 88
rect -1086 -12 -1083 -1
rect -1051 -9 -1048 -1
rect -1016 -12 -1013 -1
rect -984 -9 -981 -1
rect -953 -9 -950 -1
rect -920 -9 -917 -1
rect -1086 -14 -1013 -12
rect -1054 -87 -953 -84
rect -1089 -113 -1086 -104
rect -1054 -113 -1051 -87
rect -1019 -113 -1016 -104
rect -987 -113 -984 -104
rect -956 -113 -953 -87
rect -923 -113 -920 -104
rect -1089 -202 -1086 -119
rect -1054 -202 -1051 -119
rect -1019 -202 -1016 -119
rect -987 -202 -984 -119
rect -956 -202 -953 -119
rect -923 -202 -920 -119
rect -1089 -219 -1086 -208
rect -1054 -216 -1051 -208
rect -1019 -219 -1016 -208
rect -987 -216 -984 -208
rect -956 -216 -953 -208
rect -923 -216 -920 -208
rect -1089 -221 -1016 -219
<< polycontact >>
rect -1096 523 -1089 529
rect -1060 522 -1054 528
rect -993 522 -987 528
rect -929 498 -923 503
rect -1097 276 -1090 282
rect -1061 275 -1055 281
rect -994 275 -988 281
rect -930 251 -924 256
rect -739 208 -730 217
rect -694 207 -685 216
rect -646 206 -637 215
rect -603 206 -594 215
rect -559 204 -550 213
rect -518 212 -508 221
rect -1093 50 -1086 56
rect -1057 49 -1051 55
rect -990 49 -984 55
rect -926 25 -920 30
rect -1096 -157 -1089 -151
rect -1060 -158 -1054 -152
rect -993 -158 -987 -152
rect -929 -182 -923 -177
<< metal1 >>
rect -1117 611 -953 612
rect -1180 600 -694 611
rect -1180 365 -1173 600
rect -1099 567 -1095 600
rect -1065 567 -1061 600
rect -1032 567 -1028 600
rect -1000 567 -996 600
rect -977 599 -694 600
rect -945 586 -881 592
rect -945 567 -941 586
rect -913 567 -909 586
rect -1104 523 -1096 529
rect -1076 478 -1072 563
rect -1042 528 -1038 563
rect -1009 539 -1005 563
rect -977 539 -973 563
rect -968 539 -964 563
rect -936 539 -932 563
rect -885 542 -881 586
rect -1009 535 -932 539
rect -886 537 -769 542
rect -1067 522 -1060 528
rect -1042 522 -993 528
rect -1042 478 -1038 522
rect -933 498 -929 503
rect -885 493 -881 537
rect -977 489 -881 493
rect -977 478 -973 489
rect -913 478 -909 489
rect -1005 474 -1000 478
rect -941 474 -936 478
rect -1099 457 -1095 474
rect -1065 457 -1061 474
rect -1032 457 -1028 474
rect -968 457 -964 474
rect -1106 442 -949 457
rect -1180 354 -954 365
rect -1180 139 -1173 354
rect -1118 353 -954 354
rect -1100 320 -1096 353
rect -1066 320 -1062 353
rect -1033 320 -1029 353
rect -1001 320 -997 353
rect -946 339 -881 345
rect -946 320 -942 339
rect -914 320 -910 339
rect -1105 276 -1097 282
rect -1077 231 -1073 316
rect -1043 281 -1039 316
rect -1010 292 -1006 316
rect -978 292 -974 316
rect -969 292 -965 316
rect -937 292 -933 316
rect -1010 288 -933 292
rect -1068 275 -1061 281
rect -1043 275 -994 281
rect -1043 231 -1039 275
rect -886 268 -881 339
rect -794 268 -787 269
rect -887 263 -787 268
rect -934 251 -930 256
rect -886 246 -881 263
rect -978 242 -881 246
rect -794 243 -787 263
rect -978 231 -974 242
rect -914 231 -910 242
rect -1006 227 -1001 231
rect -942 227 -937 231
rect -1100 210 -1096 227
rect -1066 210 -1062 227
rect -1033 210 -1029 227
rect -969 211 -965 227
rect -772 216 -769 537
rect -703 301 -694 599
rect -753 292 -451 301
rect -753 286 -477 292
rect -746 274 -742 286
rect -702 274 -698 286
rect -658 274 -654 286
rect -614 274 -610 286
rect -570 274 -566 286
rect -526 274 -522 286
rect -710 259 -706 270
rect -666 259 -662 270
rect -622 259 -618 270
rect -578 259 -574 270
rect -534 259 -530 270
rect -710 255 -530 259
rect -534 221 -525 255
rect -490 224 -486 270
rect -459 246 -452 292
rect -748 216 -739 217
rect -970 210 -810 211
rect -1100 195 -810 210
rect -772 208 -739 216
rect -698 207 -694 216
rect -649 206 -646 215
rect -608 206 -603 215
rect -564 205 -559 213
rect -568 204 -559 205
rect -534 212 -518 221
rect -490 212 -478 224
rect -970 194 -810 195
rect -818 152 -810 194
rect -534 171 -530 212
rect -490 171 -486 212
rect -706 167 -702 171
rect -662 167 -658 171
rect -618 167 -614 171
rect -574 167 -570 171
rect -746 153 -742 167
rect -526 153 -522 167
rect -749 152 -473 153
rect -1180 128 -950 139
rect -818 138 -473 152
rect -1180 85 -1173 128
rect -1114 127 -950 128
rect -1096 94 -1092 127
rect -1062 94 -1058 127
rect -1029 94 -1025 127
rect -997 94 -993 127
rect -942 113 -877 119
rect -942 94 -938 113
rect -910 94 -906 113
rect -1181 -68 -1173 85
rect -1101 50 -1093 56
rect -1073 5 -1069 90
rect -1039 55 -1035 90
rect -1006 66 -1002 90
rect -974 66 -970 90
rect -882 110 -877 113
rect -882 104 -658 110
rect -965 66 -961 90
rect -933 66 -929 90
rect -1006 62 -929 66
rect -1064 49 -1057 55
rect -1039 49 -990 55
rect -1039 5 -1035 49
rect -930 25 -926 30
rect -882 20 -877 104
rect -974 16 -877 20
rect -974 5 -970 16
rect -910 5 -906 16
rect -1002 1 -997 5
rect -938 1 -933 5
rect -1096 -16 -1092 1
rect -1062 -16 -1058 1
rect -1029 -16 -1025 1
rect -965 -16 -961 1
rect -1094 -31 -946 -16
rect -1181 -79 -953 -68
rect -1117 -80 -953 -79
rect -1099 -113 -1095 -80
rect -1065 -113 -1061 -80
rect -1032 -113 -1028 -80
rect -1000 -113 -996 -80
rect -945 -94 -879 -88
rect -945 -113 -941 -94
rect -913 -113 -909 -94
rect -1104 -157 -1096 -151
rect -1076 -202 -1072 -117
rect -1042 -152 -1038 -117
rect -1009 -141 -1005 -117
rect -977 -141 -973 -117
rect -968 -141 -964 -117
rect -936 -141 -932 -117
rect -1009 -145 -932 -141
rect -885 -133 -880 -94
rect -617 -133 -605 103
rect -885 -142 -605 -133
rect -1067 -158 -1060 -152
rect -1042 -158 -993 -152
rect -1042 -202 -1038 -158
rect -933 -182 -929 -177
rect -885 -187 -880 -142
rect -977 -191 -879 -187
rect -977 -202 -973 -191
rect -913 -202 -909 -191
rect -1005 -206 -1000 -202
rect -941 -206 -936 -202
rect -1099 -222 -1095 -206
rect -1096 -223 -1095 -222
rect -1065 -223 -1061 -206
rect -1032 -223 -1028 -206
rect -968 -223 -964 -206
rect -1096 -238 -949 -223
<< m2contact >>
rect -1072 498 -1064 503
rect -940 498 -933 503
rect -1127 441 -1106 458
rect -1073 251 -1065 256
rect -941 251 -934 256
rect -794 227 -787 243
rect -1119 195 -1100 211
rect -459 232 -451 246
rect -710 207 -698 217
rect -658 205 -649 216
rect -617 205 -608 215
rect -572 205 -564 219
rect -658 104 -648 118
rect -1069 25 -1061 30
rect -937 25 -930 30
rect -618 103 -604 121
rect -1113 -32 -1094 -16
rect -1072 -182 -1064 -177
rect -940 -182 -933 -177
rect -1115 -238 -1096 -222
<< metal2 >>
rect -1064 498 -940 503
rect -1137 441 -1127 458
rect -1137 431 -1116 441
rect -1136 205 -1129 431
rect -1065 251 -941 256
rect -572 232 -459 239
rect -787 227 -703 232
rect -794 226 -703 227
rect -710 217 -703 226
rect -572 228 -451 232
rect -572 219 -564 228
rect -1136 196 -1119 205
rect -1136 -18 -1129 196
rect -658 118 -651 205
rect -614 121 -610 205
rect -1061 25 -937 30
rect -1136 -23 -1124 -18
rect -1136 -32 -1113 -23
rect -1136 -230 -1129 -32
rect -1064 -182 -940 -177
rect -1136 -238 -1115 -230
rect -1136 -239 -1111 -238
<< labels >>
rlabel metal1 -1102 524 -1102 524 1 node_a0
rlabel metal1 -1064 526 -1064 526 1 node_b0
rlabel metal1 -1102 279 -1102 279 1 node_a1
rlabel metal1 -1066 278 -1066 278 1 node_b1
rlabel metal1 -1097 52 -1097 52 1 node_a2
rlabel metal1 -1060 51 -1060 51 1 node_b2
rlabel metal1 -1102 -154 -1102 -154 1 node_a3
rlabel metal1 -1064 -155 -1064 -155 1 node_b3
rlabel metal1 -1112 604 -1112 604 1 vdd
rlabel metal1 -1027 445 -1027 445 1 gnd
rlabel metal1 -487 218 -487 218 1 node_c2
<< end >>
